module x_delay_line (
   input    logic                         i_clk,
   input    logic                         i_dl,
   input    logic [$clog2(256)-1:0]  i_sel,
   output   logic                         o_data
);

logic [256:0]   p0_dl;
logic [256-1:0] p1_dl;
logic [256-1:0] p2_dl;
logic [256-1:0] p3_dl;

assign p0_dl[0] = i_dl;

   (* BEL="X1/Y1/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut0 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[0]    ),
      .O       (p0_dl[1]  )
   );

   (* BEL="X1/Y1/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut1 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[1]    ),
      .O       (p0_dl[2]  )
   );

   (* BEL="X1/Y1/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut2 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[2]    ),
      .O       (p0_dl[3]  )
   );

   (* BEL="X1/Y1/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut3 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[3]    ),
      .O       (p0_dl[4]  )
   );

   (* BEL="X1/Y1/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut4 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[4]    ),
      .O       (p0_dl[5]  )
   );

   (* BEL="X1/Y1/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut5 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[5]    ),
      .O       (p0_dl[6]  )
   );

   (* BEL="X1/Y1/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut6 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[6]    ),
      .O       (p0_dl[7]  )
   );

   (* BEL="X1/Y1/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut7 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[7]    ),
      .O       (p0_dl[8]  )
   );

   (* BEL="X1/Y2/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut8 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[8]    ),
      .O       (p0_dl[9]  )
   );

   (* BEL="X1/Y2/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut9 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[9]    ),
      .O       (p0_dl[10]  )
   );

   (* BEL="X1/Y2/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut10 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[10]    ),
      .O       (p0_dl[11]  )
   );

   (* BEL="X1/Y2/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut11 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[11]    ),
      .O       (p0_dl[12]  )
   );

   (* BEL="X1/Y2/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut12 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[12]    ),
      .O       (p0_dl[13]  )
   );

   (* BEL="X1/Y2/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut13 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[13]    ),
      .O       (p0_dl[14]  )
   );

   (* BEL="X1/Y2/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut14 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[14]    ),
      .O       (p0_dl[15]  )
   );

   (* BEL="X1/Y2/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut15 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[15]    ),
      .O       (p0_dl[16]  )
   );

   (* BEL="X1/Y3/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut16 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[16]    ),
      .O       (p0_dl[17]  )
   );

   (* BEL="X1/Y3/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut17 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[17]    ),
      .O       (p0_dl[18]  )
   );

   (* BEL="X1/Y3/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut18 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[18]    ),
      .O       (p0_dl[19]  )
   );

   (* BEL="X1/Y3/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut19 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[19]    ),
      .O       (p0_dl[20]  )
   );

   (* BEL="X1/Y3/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut20 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[20]    ),
      .O       (p0_dl[21]  )
   );

   (* BEL="X1/Y3/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut21 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[21]    ),
      .O       (p0_dl[22]  )
   );

   (* BEL="X1/Y3/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut22 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[22]    ),
      .O       (p0_dl[23]  )
   );

   (* BEL="X1/Y3/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut23 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[23]    ),
      .O       (p0_dl[24]  )
   );

   (* BEL="X1/Y4/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut24 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[24]    ),
      .O       (p0_dl[25]  )
   );

   (* BEL="X1/Y4/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut25 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[25]    ),
      .O       (p0_dl[26]  )
   );

   (* BEL="X1/Y4/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut26 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[26]    ),
      .O       (p0_dl[27]  )
   );

   (* BEL="X1/Y4/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut27 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[27]    ),
      .O       (p0_dl[28]  )
   );

   (* BEL="X1/Y4/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut28 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[28]    ),
      .O       (p0_dl[29]  )
   );

   (* BEL="X1/Y4/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut29 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[29]    ),
      .O       (p0_dl[30]  )
   );

   (* BEL="X1/Y4/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut30 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[30]    ),
      .O       (p0_dl[31]  )
   );

   (* BEL="X1/Y4/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut31 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[31]    ),
      .O       (p0_dl[32]  )
   );

   (* BEL="X1/Y5/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut32 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[32]    ),
      .O       (p0_dl[33]  )
   );

   (* BEL="X1/Y5/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut33 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[33]    ),
      .O       (p0_dl[34]  )
   );

   (* BEL="X1/Y5/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut34 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[34]    ),
      .O       (p0_dl[35]  )
   );

   (* BEL="X1/Y5/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut35 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[35]    ),
      .O       (p0_dl[36]  )
   );

   (* BEL="X1/Y5/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut36 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[36]    ),
      .O       (p0_dl[37]  )
   );

   (* BEL="X1/Y5/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut37 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[37]    ),
      .O       (p0_dl[38]  )
   );

   (* BEL="X1/Y5/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut38 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[38]    ),
      .O       (p0_dl[39]  )
   );

   (* BEL="X1/Y5/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut39 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[39]    ),
      .O       (p0_dl[40]  )
   );

   (* BEL="X1/Y6/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut40 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[40]    ),
      .O       (p0_dl[41]  )
   );

   (* BEL="X1/Y6/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut41 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[41]    ),
      .O       (p0_dl[42]  )
   );

   (* BEL="X1/Y6/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut42 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[42]    ),
      .O       (p0_dl[43]  )
   );

   (* BEL="X1/Y6/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut43 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[43]    ),
      .O       (p0_dl[44]  )
   );

   (* BEL="X1/Y6/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut44 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[44]    ),
      .O       (p0_dl[45]  )
   );

   (* BEL="X1/Y6/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut45 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[45]    ),
      .O       (p0_dl[46]  )
   );

   (* BEL="X1/Y6/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut46 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[46]    ),
      .O       (p0_dl[47]  )
   );

   (* BEL="X1/Y6/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut47 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[47]    ),
      .O       (p0_dl[48]  )
   );

   (* BEL="X1/Y7/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut48 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[48]    ),
      .O       (p0_dl[49]  )
   );

   (* BEL="X1/Y7/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut49 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[49]    ),
      .O       (p0_dl[50]  )
   );

   (* BEL="X1/Y7/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut50 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[50]    ),
      .O       (p0_dl[51]  )
   );

   (* BEL="X1/Y7/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut51 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[51]    ),
      .O       (p0_dl[52]  )
   );

   (* BEL="X1/Y7/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut52 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[52]    ),
      .O       (p0_dl[53]  )
   );

   (* BEL="X1/Y7/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut53 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[53]    ),
      .O       (p0_dl[54]  )
   );

   (* BEL="X1/Y7/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut54 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[54]    ),
      .O       (p0_dl[55]  )
   );

   (* BEL="X1/Y7/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut55 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[55]    ),
      .O       (p0_dl[56]  )
   );

   (* BEL="X1/Y8/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut56 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[56]    ),
      .O       (p0_dl[57]  )
   );

   (* BEL="X1/Y8/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut57 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[57]    ),
      .O       (p0_dl[58]  )
   );

   (* BEL="X1/Y8/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut58 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[58]    ),
      .O       (p0_dl[59]  )
   );

   (* BEL="X1/Y8/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut59 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[59]    ),
      .O       (p0_dl[60]  )
   );

   (* BEL="X1/Y8/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut60 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[60]    ),
      .O       (p0_dl[61]  )
   );

   (* BEL="X1/Y8/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut61 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[61]    ),
      .O       (p0_dl[62]  )
   );

   (* BEL="X1/Y8/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut62 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[62]    ),
      .O       (p0_dl[63]  )
   );

   (* BEL="X1/Y8/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut63 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[63]    ),
      .O       (p0_dl[64]  )
   );

   (* BEL="X1/Y9/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut64 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[64]    ),
      .O       (p0_dl[65]  )
   );

   (* BEL="X1/Y9/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut65 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[65]    ),
      .O       (p0_dl[66]  )
   );

   (* BEL="X1/Y9/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut66 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[66]    ),
      .O       (p0_dl[67]  )
   );

   (* BEL="X1/Y9/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut67 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[67]    ),
      .O       (p0_dl[68]  )
   );

   (* BEL="X1/Y9/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut68 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[68]    ),
      .O       (p0_dl[69]  )
   );

   (* BEL="X1/Y9/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut69 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[69]    ),
      .O       (p0_dl[70]  )
   );

   (* BEL="X1/Y9/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut70 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[70]    ),
      .O       (p0_dl[71]  )
   );

   (* BEL="X1/Y9/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut71 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[71]    ),
      .O       (p0_dl[72]  )
   );

   (* BEL="X1/Y10/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut72 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[72]    ),
      .O       (p0_dl[73]  )
   );

   (* BEL="X1/Y10/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut73 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[73]    ),
      .O       (p0_dl[74]  )
   );

   (* BEL="X1/Y10/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut74 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[74]    ),
      .O       (p0_dl[75]  )
   );

   (* BEL="X1/Y10/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut75 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[75]    ),
      .O       (p0_dl[76]  )
   );

   (* BEL="X1/Y10/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut76 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[76]    ),
      .O       (p0_dl[77]  )
   );

   (* BEL="X1/Y10/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut77 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[77]    ),
      .O       (p0_dl[78]  )
   );

   (* BEL="X1/Y10/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut78 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[78]    ),
      .O       (p0_dl[79]  )
   );

   (* BEL="X1/Y10/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut79 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[79]    ),
      .O       (p0_dl[80]  )
   );

   (* BEL="X1/Y11/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut80 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[80]    ),
      .O       (p0_dl[81]  )
   );

   (* BEL="X1/Y11/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut81 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[81]    ),
      .O       (p0_dl[82]  )
   );

   (* BEL="X1/Y11/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut82 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[82]    ),
      .O       (p0_dl[83]  )
   );

   (* BEL="X1/Y11/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut83 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[83]    ),
      .O       (p0_dl[84]  )
   );

   (* BEL="X1/Y11/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut84 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[84]    ),
      .O       (p0_dl[85]  )
   );

   (* BEL="X1/Y11/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut85 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[85]    ),
      .O       (p0_dl[86]  )
   );

   (* BEL="X1/Y11/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut86 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[86]    ),
      .O       (p0_dl[87]  )
   );

   (* BEL="X1/Y11/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut87 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[87]    ),
      .O       (p0_dl[88]  )
   );

   (* BEL="X1/Y12/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut88 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[88]    ),
      .O       (p0_dl[89]  )
   );

   (* BEL="X1/Y12/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut89 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[89]    ),
      .O       (p0_dl[90]  )
   );

   (* BEL="X1/Y12/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut90 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[90]    ),
      .O       (p0_dl[91]  )
   );

   (* BEL="X1/Y12/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut91 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[91]    ),
      .O       (p0_dl[92]  )
   );

   (* BEL="X1/Y12/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut92 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[92]    ),
      .O       (p0_dl[93]  )
   );

   (* BEL="X1/Y12/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut93 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[93]    ),
      .O       (p0_dl[94]  )
   );

   (* BEL="X1/Y12/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut94 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[94]    ),
      .O       (p0_dl[95]  )
   );

   (* BEL="X1/Y12/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut95 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[95]    ),
      .O       (p0_dl[96]  )
   );

   (* BEL="X1/Y13/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut96 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[96]    ),
      .O       (p0_dl[97]  )
   );

   (* BEL="X1/Y13/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut97 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[97]    ),
      .O       (p0_dl[98]  )
   );

   (* BEL="X1/Y13/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut98 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[98]    ),
      .O       (p0_dl[99]  )
   );

   (* BEL="X1/Y13/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut99 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[99]    ),
      .O       (p0_dl[100]  )
   );

   (* BEL="X1/Y13/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut100 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[100]    ),
      .O       (p0_dl[101]  )
   );

   (* BEL="X1/Y13/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut101 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[101]    ),
      .O       (p0_dl[102]  )
   );

   (* BEL="X1/Y13/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut102 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[102]    ),
      .O       (p0_dl[103]  )
   );

   (* BEL="X1/Y13/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut103 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[103]    ),
      .O       (p0_dl[104]  )
   );

   (* BEL="X1/Y14/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut104 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[104]    ),
      .O       (p0_dl[105]  )
   );

   (* BEL="X1/Y14/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut105 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[105]    ),
      .O       (p0_dl[106]  )
   );

   (* BEL="X1/Y14/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut106 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[106]    ),
      .O       (p0_dl[107]  )
   );

   (* BEL="X1/Y14/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut107 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[107]    ),
      .O       (p0_dl[108]  )
   );

   (* BEL="X1/Y14/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut108 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[108]    ),
      .O       (p0_dl[109]  )
   );

   (* BEL="X1/Y14/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut109 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[109]    ),
      .O       (p0_dl[110]  )
   );

   (* BEL="X1/Y14/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut110 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[110]    ),
      .O       (p0_dl[111]  )
   );

   (* BEL="X1/Y14/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut111 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[111]    ),
      .O       (p0_dl[112]  )
   );

   (* BEL="X1/Y15/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut112 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[112]    ),
      .O       (p0_dl[113]  )
   );

   (* BEL="X1/Y15/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut113 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[113]    ),
      .O       (p0_dl[114]  )
   );

   (* BEL="X1/Y15/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut114 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[114]    ),
      .O       (p0_dl[115]  )
   );

   (* BEL="X1/Y15/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut115 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[115]    ),
      .O       (p0_dl[116]  )
   );

   (* BEL="X1/Y15/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut116 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[116]    ),
      .O       (p0_dl[117]  )
   );

   (* BEL="X1/Y15/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut117 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[117]    ),
      .O       (p0_dl[118]  )
   );

   (* BEL="X1/Y15/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut118 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[118]    ),
      .O       (p0_dl[119]  )
   );

   (* BEL="X1/Y15/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut119 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[119]    ),
      .O       (p0_dl[120]  )
   );

   (* BEL="X1/Y16/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut120 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[120]    ),
      .O       (p0_dl[121]  )
   );

   (* BEL="X1/Y16/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut121 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[121]    ),
      .O       (p0_dl[122]  )
   );

   (* BEL="X1/Y16/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut122 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[122]    ),
      .O       (p0_dl[123]  )
   );

   (* BEL="X1/Y16/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut123 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[123]    ),
      .O       (p0_dl[124]  )
   );

   (* BEL="X1/Y16/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut124 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[124]    ),
      .O       (p0_dl[125]  )
   );

   (* BEL="X1/Y16/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut125 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[125]    ),
      .O       (p0_dl[126]  )
   );

   (* BEL="X1/Y16/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut126 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[126]    ),
      .O       (p0_dl[127]  )
   );

   (* BEL="X1/Y16/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut127 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[127]    ),
      .O       (p0_dl[128]  )
   );

   (* BEL="X1/Y17/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut128 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[128]    ),
      .O       (p0_dl[129]  )
   );

   (* BEL="X1/Y17/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut129 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[129]    ),
      .O       (p0_dl[130]  )
   );

   (* BEL="X1/Y17/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut130 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[130]    ),
      .O       (p0_dl[131]  )
   );

   (* BEL="X1/Y17/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut131 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[131]    ),
      .O       (p0_dl[132]  )
   );

   (* BEL="X1/Y17/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut132 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[132]    ),
      .O       (p0_dl[133]  )
   );

   (* BEL="X1/Y17/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut133 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[133]    ),
      .O       (p0_dl[134]  )
   );

   (* BEL="X1/Y17/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut134 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[134]    ),
      .O       (p0_dl[135]  )
   );

   (* BEL="X1/Y17/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut135 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[135]    ),
      .O       (p0_dl[136]  )
   );

   (* BEL="X1/Y18/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut136 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[136]    ),
      .O       (p0_dl[137]  )
   );

   (* BEL="X1/Y18/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut137 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[137]    ),
      .O       (p0_dl[138]  )
   );

   (* BEL="X1/Y18/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut138 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[138]    ),
      .O       (p0_dl[139]  )
   );

   (* BEL="X1/Y18/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut139 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[139]    ),
      .O       (p0_dl[140]  )
   );

   (* BEL="X1/Y18/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut140 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[140]    ),
      .O       (p0_dl[141]  )
   );

   (* BEL="X1/Y18/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut141 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[141]    ),
      .O       (p0_dl[142]  )
   );

   (* BEL="X1/Y18/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut142 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[142]    ),
      .O       (p0_dl[143]  )
   );

   (* BEL="X1/Y18/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut143 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[143]    ),
      .O       (p0_dl[144]  )
   );

   (* BEL="X1/Y19/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut144 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[144]    ),
      .O       (p0_dl[145]  )
   );

   (* BEL="X1/Y19/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut145 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[145]    ),
      .O       (p0_dl[146]  )
   );

   (* BEL="X1/Y19/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut146 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[146]    ),
      .O       (p0_dl[147]  )
   );

   (* BEL="X1/Y19/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut147 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[147]    ),
      .O       (p0_dl[148]  )
   );

   (* BEL="X1/Y19/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut148 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[148]    ),
      .O       (p0_dl[149]  )
   );

   (* BEL="X1/Y19/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut149 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[149]    ),
      .O       (p0_dl[150]  )
   );

   (* BEL="X1/Y19/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut150 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[150]    ),
      .O       (p0_dl[151]  )
   );

   (* BEL="X1/Y19/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut151 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[151]    ),
      .O       (p0_dl[152]  )
   );

   (* BEL="X1/Y20/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut152 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[152]    ),
      .O       (p0_dl[153]  )
   );

   (* BEL="X1/Y20/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut153 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[153]    ),
      .O       (p0_dl[154]  )
   );

   (* BEL="X1/Y20/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut154 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[154]    ),
      .O       (p0_dl[155]  )
   );

   (* BEL="X1/Y20/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut155 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[155]    ),
      .O       (p0_dl[156]  )
   );

   (* BEL="X1/Y20/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut156 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[156]    ),
      .O       (p0_dl[157]  )
   );

   (* BEL="X1/Y20/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut157 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[157]    ),
      .O       (p0_dl[158]  )
   );

   (* BEL="X1/Y20/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut158 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[158]    ),
      .O       (p0_dl[159]  )
   );

   (* BEL="X1/Y20/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut159 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[159]    ),
      .O       (p0_dl[160]  )
   );

   (* BEL="X1/Y21/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut160 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[160]    ),
      .O       (p0_dl[161]  )
   );

   (* BEL="X1/Y21/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut161 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[161]    ),
      .O       (p0_dl[162]  )
   );

   (* BEL="X1/Y21/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut162 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[162]    ),
      .O       (p0_dl[163]  )
   );

   (* BEL="X1/Y21/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut163 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[163]    ),
      .O       (p0_dl[164]  )
   );

   (* BEL="X1/Y21/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut164 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[164]    ),
      .O       (p0_dl[165]  )
   );

   (* BEL="X1/Y21/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut165 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[165]    ),
      .O       (p0_dl[166]  )
   );

   (* BEL="X1/Y21/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut166 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[166]    ),
      .O       (p0_dl[167]  )
   );

   (* BEL="X1/Y21/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut167 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[167]    ),
      .O       (p0_dl[168]  )
   );

   (* BEL="X1/Y22/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut168 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[168]    ),
      .O       (p0_dl[169]  )
   );

   (* BEL="X1/Y22/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut169 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[169]    ),
      .O       (p0_dl[170]  )
   );

   (* BEL="X1/Y22/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut170 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[170]    ),
      .O       (p0_dl[171]  )
   );

   (* BEL="X1/Y22/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut171 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[171]    ),
      .O       (p0_dl[172]  )
   );

   (* BEL="X1/Y22/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut172 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[172]    ),
      .O       (p0_dl[173]  )
   );

   (* BEL="X1/Y22/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut173 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[173]    ),
      .O       (p0_dl[174]  )
   );

   (* BEL="X1/Y22/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut174 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[174]    ),
      .O       (p0_dl[175]  )
   );

   (* BEL="X1/Y22/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut175 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[175]    ),
      .O       (p0_dl[176]  )
   );

   (* BEL="X1/Y23/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut176 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[176]    ),
      .O       (p0_dl[177]  )
   );

   (* BEL="X1/Y23/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut177 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[177]    ),
      .O       (p0_dl[178]  )
   );

   (* BEL="X1/Y23/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut178 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[178]    ),
      .O       (p0_dl[179]  )
   );

   (* BEL="X1/Y23/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut179 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[179]    ),
      .O       (p0_dl[180]  )
   );

   (* BEL="X1/Y23/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut180 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[180]    ),
      .O       (p0_dl[181]  )
   );

   (* BEL="X1/Y23/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut181 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[181]    ),
      .O       (p0_dl[182]  )
   );

   (* BEL="X1/Y23/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut182 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[182]    ),
      .O       (p0_dl[183]  )
   );

   (* BEL="X1/Y23/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut183 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[183]    ),
      .O       (p0_dl[184]  )
   );

   (* BEL="X1/Y24/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut184 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[184]    ),
      .O       (p0_dl[185]  )
   );

   (* BEL="X1/Y24/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut185 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[185]    ),
      .O       (p0_dl[186]  )
   );

   (* BEL="X1/Y24/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut186 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[186]    ),
      .O       (p0_dl[187]  )
   );

   (* BEL="X1/Y24/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut187 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[187]    ),
      .O       (p0_dl[188]  )
   );

   (* BEL="X1/Y24/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut188 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[188]    ),
      .O       (p0_dl[189]  )
   );

   (* BEL="X1/Y24/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut189 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[189]    ),
      .O       (p0_dl[190]  )
   );

   (* BEL="X1/Y24/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut190 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[190]    ),
      .O       (p0_dl[191]  )
   );

   (* BEL="X1/Y24/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut191 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[191]    ),
      .O       (p0_dl[192]  )
   );

   (* BEL="X1/Y25/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut192 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[192]    ),
      .O       (p0_dl[193]  )
   );

   (* BEL="X1/Y25/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut193 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[193]    ),
      .O       (p0_dl[194]  )
   );

   (* BEL="X1/Y25/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut194 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[194]    ),
      .O       (p0_dl[195]  )
   );

   (* BEL="X1/Y25/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut195 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[195]    ),
      .O       (p0_dl[196]  )
   );

   (* BEL="X1/Y25/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut196 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[196]    ),
      .O       (p0_dl[197]  )
   );

   (* BEL="X1/Y25/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut197 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[197]    ),
      .O       (p0_dl[198]  )
   );

   (* BEL="X1/Y25/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut198 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[198]    ),
      .O       (p0_dl[199]  )
   );

   (* BEL="X1/Y25/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut199 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[199]    ),
      .O       (p0_dl[200]  )
   );

   (* BEL="X1/Y26/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut200 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[200]    ),
      .O       (p0_dl[201]  )
   );

   (* BEL="X1/Y26/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut201 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[201]    ),
      .O       (p0_dl[202]  )
   );

   (* BEL="X1/Y26/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut202 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[202]    ),
      .O       (p0_dl[203]  )
   );

   (* BEL="X1/Y26/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut203 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[203]    ),
      .O       (p0_dl[204]  )
   );

   (* BEL="X1/Y26/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut204 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[204]    ),
      .O       (p0_dl[205]  )
   );

   (* BEL="X1/Y26/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut205 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[205]    ),
      .O       (p0_dl[206]  )
   );

   (* BEL="X1/Y26/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut206 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[206]    ),
      .O       (p0_dl[207]  )
   );

   (* BEL="X1/Y26/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut207 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[207]    ),
      .O       (p0_dl[208]  )
   );

   (* BEL="X1/Y27/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut208 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[208]    ),
      .O       (p0_dl[209]  )
   );

   (* BEL="X1/Y27/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut209 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[209]    ),
      .O       (p0_dl[210]  )
   );

   (* BEL="X1/Y27/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut210 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[210]    ),
      .O       (p0_dl[211]  )
   );

   (* BEL="X1/Y27/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut211 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[211]    ),
      .O       (p0_dl[212]  )
   );

   (* BEL="X1/Y27/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut212 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[212]    ),
      .O       (p0_dl[213]  )
   );

   (* BEL="X1/Y27/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut213 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[213]    ),
      .O       (p0_dl[214]  )
   );

   (* BEL="X1/Y27/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut214 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[214]    ),
      .O       (p0_dl[215]  )
   );

   (* BEL="X1/Y27/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut215 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[215]    ),
      .O       (p0_dl[216]  )
   );

   (* BEL="X1/Y28/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut216 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[216]    ),
      .O       (p0_dl[217]  )
   );

   (* BEL="X1/Y28/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut217 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[217]    ),
      .O       (p0_dl[218]  )
   );

   (* BEL="X1/Y28/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut218 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[218]    ),
      .O       (p0_dl[219]  )
   );

   (* BEL="X1/Y28/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut219 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[219]    ),
      .O       (p0_dl[220]  )
   );

   (* BEL="X1/Y28/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut220 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[220]    ),
      .O       (p0_dl[221]  )
   );

   (* BEL="X1/Y28/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut221 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[221]    ),
      .O       (p0_dl[222]  )
   );

   (* BEL="X1/Y28/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut222 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[222]    ),
      .O       (p0_dl[223]  )
   );

   (* BEL="X1/Y28/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut223 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[223]    ),
      .O       (p0_dl[224]  )
   );

   (* BEL="X1/Y29/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut224 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[224]    ),
      .O       (p0_dl[225]  )
   );

   (* BEL="X1/Y29/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut225 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[225]    ),
      .O       (p0_dl[226]  )
   );

   (* BEL="X1/Y29/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut226 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[226]    ),
      .O       (p0_dl[227]  )
   );

   (* BEL="X1/Y29/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut227 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[227]    ),
      .O       (p0_dl[228]  )
   );

   (* BEL="X1/Y29/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut228 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[228]    ),
      .O       (p0_dl[229]  )
   );

   (* BEL="X1/Y29/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut229 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[229]    ),
      .O       (p0_dl[230]  )
   );

   (* BEL="X1/Y29/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut230 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[230]    ),
      .O       (p0_dl[231]  )
   );

   (* BEL="X1/Y29/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut231 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[231]    ),
      .O       (p0_dl[232]  )
   );

   (* BEL="X1/Y30/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut232 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[232]    ),
      .O       (p0_dl[233]  )
   );

   (* BEL="X1/Y30/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut233 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[233]    ),
      .O       (p0_dl[234]  )
   );

   (* BEL="X1/Y30/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut234 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[234]    ),
      .O       (p0_dl[235]  )
   );

   (* BEL="X1/Y30/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut235 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[235]    ),
      .O       (p0_dl[236]  )
   );

   (* BEL="X1/Y30/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut236 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[236]    ),
      .O       (p0_dl[237]  )
   );

   (* BEL="X1/Y30/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut237 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[237]    ),
      .O       (p0_dl[238]  )
   );

   (* BEL="X1/Y30/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut238 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[238]    ),
      .O       (p0_dl[239]  )
   );

   (* BEL="X1/Y30/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut239 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[239]    ),
      .O       (p0_dl[240]  )
   );

   (* BEL="X1/Y31/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut240 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[240]    ),
      .O       (p0_dl[241]  )
   );

   (* BEL="X1/Y31/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut241 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[241]    ),
      .O       (p0_dl[242]  )
   );

   (* BEL="X1/Y31/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut242 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[242]    ),
      .O       (p0_dl[243]  )
   );

   (* BEL="X1/Y31/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut243 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[243]    ),
      .O       (p0_dl[244]  )
   );

   (* BEL="X1/Y31/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut244 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[244]    ),
      .O       (p0_dl[245]  )
   );

   (* BEL="X1/Y31/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut245 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[245]    ),
      .O       (p0_dl[246]  )
   );

   (* BEL="X1/Y31/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut246 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[246]    ),
      .O       (p0_dl[247]  )
   );

   (* BEL="X1/Y31/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut247 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[247]    ),
      .O       (p0_dl[248]  )
   );

   (* BEL="X1/Y32/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut248 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[248]    ),
      .O       (p0_dl[249]  )
   );

   (* BEL="X1/Y32/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut249 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[249]    ),
      .O       (p0_dl[250]  )
   );

   (* BEL="X1/Y32/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut250 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[250]    ),
      .O       (p0_dl[251]  )
   );

   (* BEL="X1/Y32/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut251 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[251]    ),
      .O       (p0_dl[252]  )
   );

   (* BEL="X1/Y32/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut252 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[252]    ),
      .O       (p0_dl[253]  )
   );

   (* BEL="X1/Y32/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut253 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[253]    ),
      .O       (p0_dl[254]  )
   );

   (* BEL="X1/Y32/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut254 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[254]    ),
      .O       (p0_dl[255]  )
   );

   (* BEL="X1/Y32/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0001      )
   ) lut255 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[255]    ),
      .O       (p0_dl[256]  )
   );


   (* BEL="X2/Y1/lc0" *)
   SB_DFF  dff_2_0 (
      .C       (i_clk         ),
      .D       (p0_dl[1]  ),
      .Q       (p1_dl[0]    )
   );

   (* BEL="X3/Y1/lc0" *)
   SB_DFF  dff_3_0 (
      .C       (i_clk         ),
      .D       (p1_dl[0]    ),
      .Q       (p2_dl[0]    )
   );


   (* BEL="X29/Y1/lc0" *)
   SB_DFF  dff_29_0 (
      .C       (i_clk         ),
      .D       (p2_dl[0]    ),
      .Q       (p3_dl[0]    )
   );
   (* BEL="X2/Y1/lc1" *)
   SB_DFF  dff_2_1 (
      .C       (i_clk         ),
      .D       (p0_dl[2]  ),
      .Q       (p1_dl[1]    )
   );

   (* BEL="X3/Y1/lc1" *)
   SB_DFF  dff_3_1 (
      .C       (i_clk         ),
      .D       (p1_dl[1]    ),
      .Q       (p2_dl[1]    )
   );


   (* BEL="X29/Y1/lc1" *)
   SB_DFF  dff_29_1 (
      .C       (i_clk         ),
      .D       (p2_dl[1]    ),
      .Q       (p3_dl[1]    )
   );
   (* BEL="X2/Y1/lc2" *)
   SB_DFF  dff_2_2 (
      .C       (i_clk         ),
      .D       (p0_dl[3]  ),
      .Q       (p1_dl[2]    )
   );

   (* BEL="X3/Y1/lc2" *)
   SB_DFF  dff_3_2 (
      .C       (i_clk         ),
      .D       (p1_dl[2]    ),
      .Q       (p2_dl[2]    )
   );


   (* BEL="X29/Y1/lc2" *)
   SB_DFF  dff_29_2 (
      .C       (i_clk         ),
      .D       (p2_dl[2]    ),
      .Q       (p3_dl[2]    )
   );
   (* BEL="X2/Y1/lc3" *)
   SB_DFF  dff_2_3 (
      .C       (i_clk         ),
      .D       (p0_dl[4]  ),
      .Q       (p1_dl[3]    )
   );

   (* BEL="X3/Y1/lc3" *)
   SB_DFF  dff_3_3 (
      .C       (i_clk         ),
      .D       (p1_dl[3]    ),
      .Q       (p2_dl[3]    )
   );


   (* BEL="X29/Y1/lc3" *)
   SB_DFF  dff_29_3 (
      .C       (i_clk         ),
      .D       (p2_dl[3]    ),
      .Q       (p3_dl[3]    )
   );
   (* BEL="X2/Y1/lc4" *)
   SB_DFF  dff_2_4 (
      .C       (i_clk         ),
      .D       (p0_dl[5]  ),
      .Q       (p1_dl[4]    )
   );

   (* BEL="X3/Y1/lc4" *)
   SB_DFF  dff_3_4 (
      .C       (i_clk         ),
      .D       (p1_dl[4]    ),
      .Q       (p2_dl[4]    )
   );


   (* BEL="X29/Y1/lc4" *)
   SB_DFF  dff_29_4 (
      .C       (i_clk         ),
      .D       (p2_dl[4]    ),
      .Q       (p3_dl[4]    )
   );
   (* BEL="X2/Y1/lc5" *)
   SB_DFF  dff_2_5 (
      .C       (i_clk         ),
      .D       (p0_dl[6]  ),
      .Q       (p1_dl[5]    )
   );

   (* BEL="X3/Y1/lc5" *)
   SB_DFF  dff_3_5 (
      .C       (i_clk         ),
      .D       (p1_dl[5]    ),
      .Q       (p2_dl[5]    )
   );


   (* BEL="X29/Y1/lc5" *)
   SB_DFF  dff_29_5 (
      .C       (i_clk         ),
      .D       (p2_dl[5]    ),
      .Q       (p3_dl[5]    )
   );
   (* BEL="X2/Y1/lc6" *)
   SB_DFF  dff_2_6 (
      .C       (i_clk         ),
      .D       (p0_dl[7]  ),
      .Q       (p1_dl[6]    )
   );

   (* BEL="X3/Y1/lc6" *)
   SB_DFF  dff_3_6 (
      .C       (i_clk         ),
      .D       (p1_dl[6]    ),
      .Q       (p2_dl[6]    )
   );


   (* BEL="X29/Y1/lc6" *)
   SB_DFF  dff_29_6 (
      .C       (i_clk         ),
      .D       (p2_dl[6]    ),
      .Q       (p3_dl[6]    )
   );
   (* BEL="X2/Y1/lc7" *)
   SB_DFF  dff_2_7 (
      .C       (i_clk         ),
      .D       (p0_dl[8]  ),
      .Q       (p1_dl[7]    )
   );

   (* BEL="X3/Y1/lc7" *)
   SB_DFF  dff_3_7 (
      .C       (i_clk         ),
      .D       (p1_dl[7]    ),
      .Q       (p2_dl[7]    )
   );


   (* BEL="X29/Y1/lc7" *)
   SB_DFF  dff_29_7 (
      .C       (i_clk         ),
      .D       (p2_dl[7]    ),
      .Q       (p3_dl[7]    )
   );
   (* BEL="X2/Y2/lc0" *)
   SB_DFF  dff_2_8 (
      .C       (i_clk         ),
      .D       (p0_dl[9]  ),
      .Q       (p1_dl[8]    )
   );

   (* BEL="X3/Y2/lc0" *)
   SB_DFF  dff_3_8 (
      .C       (i_clk         ),
      .D       (p1_dl[8]    ),
      .Q       (p2_dl[8]    )
   );


   (* BEL="X29/Y2/lc0" *)
   SB_DFF  dff_29_8 (
      .C       (i_clk         ),
      .D       (p2_dl[8]    ),
      .Q       (p3_dl[8]    )
   );
   (* BEL="X2/Y2/lc1" *)
   SB_DFF  dff_2_9 (
      .C       (i_clk         ),
      .D       (p0_dl[10]  ),
      .Q       (p1_dl[9]    )
   );

   (* BEL="X3/Y2/lc1" *)
   SB_DFF  dff_3_9 (
      .C       (i_clk         ),
      .D       (p1_dl[9]    ),
      .Q       (p2_dl[9]    )
   );


   (* BEL="X29/Y2/lc1" *)
   SB_DFF  dff_29_9 (
      .C       (i_clk         ),
      .D       (p2_dl[9]    ),
      .Q       (p3_dl[9]    )
   );
   (* BEL="X2/Y2/lc2" *)
   SB_DFF  dff_2_10 (
      .C       (i_clk         ),
      .D       (p0_dl[11]  ),
      .Q       (p1_dl[10]    )
   );

   (* BEL="X3/Y2/lc2" *)
   SB_DFF  dff_3_10 (
      .C       (i_clk         ),
      .D       (p1_dl[10]    ),
      .Q       (p2_dl[10]    )
   );


   (* BEL="X29/Y2/lc2" *)
   SB_DFF  dff_29_10 (
      .C       (i_clk         ),
      .D       (p2_dl[10]    ),
      .Q       (p3_dl[10]    )
   );
   (* BEL="X2/Y2/lc3" *)
   SB_DFF  dff_2_11 (
      .C       (i_clk         ),
      .D       (p0_dl[12]  ),
      .Q       (p1_dl[11]    )
   );

   (* BEL="X3/Y2/lc3" *)
   SB_DFF  dff_3_11 (
      .C       (i_clk         ),
      .D       (p1_dl[11]    ),
      .Q       (p2_dl[11]    )
   );


   (* BEL="X29/Y2/lc3" *)
   SB_DFF  dff_29_11 (
      .C       (i_clk         ),
      .D       (p2_dl[11]    ),
      .Q       (p3_dl[11]    )
   );
   (* BEL="X2/Y2/lc4" *)
   SB_DFF  dff_2_12 (
      .C       (i_clk         ),
      .D       (p0_dl[13]  ),
      .Q       (p1_dl[12]    )
   );

   (* BEL="X3/Y2/lc4" *)
   SB_DFF  dff_3_12 (
      .C       (i_clk         ),
      .D       (p1_dl[12]    ),
      .Q       (p2_dl[12]    )
   );


   (* BEL="X29/Y2/lc4" *)
   SB_DFF  dff_29_12 (
      .C       (i_clk         ),
      .D       (p2_dl[12]    ),
      .Q       (p3_dl[12]    )
   );
   (* BEL="X2/Y2/lc5" *)
   SB_DFF  dff_2_13 (
      .C       (i_clk         ),
      .D       (p0_dl[14]  ),
      .Q       (p1_dl[13]    )
   );

   (* BEL="X3/Y2/lc5" *)
   SB_DFF  dff_3_13 (
      .C       (i_clk         ),
      .D       (p1_dl[13]    ),
      .Q       (p2_dl[13]    )
   );


   (* BEL="X29/Y2/lc5" *)
   SB_DFF  dff_29_13 (
      .C       (i_clk         ),
      .D       (p2_dl[13]    ),
      .Q       (p3_dl[13]    )
   );
   (* BEL="X2/Y2/lc6" *)
   SB_DFF  dff_2_14 (
      .C       (i_clk         ),
      .D       (p0_dl[15]  ),
      .Q       (p1_dl[14]    )
   );

   (* BEL="X3/Y2/lc6" *)
   SB_DFF  dff_3_14 (
      .C       (i_clk         ),
      .D       (p1_dl[14]    ),
      .Q       (p2_dl[14]    )
   );


   (* BEL="X29/Y2/lc6" *)
   SB_DFF  dff_29_14 (
      .C       (i_clk         ),
      .D       (p2_dl[14]    ),
      .Q       (p3_dl[14]    )
   );
   (* BEL="X2/Y2/lc7" *)
   SB_DFF  dff_2_15 (
      .C       (i_clk         ),
      .D       (p0_dl[16]  ),
      .Q       (p1_dl[15]    )
   );

   (* BEL="X3/Y2/lc7" *)
   SB_DFF  dff_3_15 (
      .C       (i_clk         ),
      .D       (p1_dl[15]    ),
      .Q       (p2_dl[15]    )
   );


   (* BEL="X29/Y2/lc7" *)
   SB_DFF  dff_29_15 (
      .C       (i_clk         ),
      .D       (p2_dl[15]    ),
      .Q       (p3_dl[15]    )
   );
   (* BEL="X2/Y3/lc0" *)
   SB_DFF  dff_2_16 (
      .C       (i_clk         ),
      .D       (p0_dl[17]  ),
      .Q       (p1_dl[16]    )
   );

   (* BEL="X3/Y3/lc0" *)
   SB_DFF  dff_3_16 (
      .C       (i_clk         ),
      .D       (p1_dl[16]    ),
      .Q       (p2_dl[16]    )
   );


   (* BEL="X29/Y3/lc0" *)
   SB_DFF  dff_29_16 (
      .C       (i_clk         ),
      .D       (p2_dl[16]    ),
      .Q       (p3_dl[16]    )
   );
   (* BEL="X2/Y3/lc1" *)
   SB_DFF  dff_2_17 (
      .C       (i_clk         ),
      .D       (p0_dl[18]  ),
      .Q       (p1_dl[17]    )
   );

   (* BEL="X3/Y3/lc1" *)
   SB_DFF  dff_3_17 (
      .C       (i_clk         ),
      .D       (p1_dl[17]    ),
      .Q       (p2_dl[17]    )
   );


   (* BEL="X29/Y3/lc1" *)
   SB_DFF  dff_29_17 (
      .C       (i_clk         ),
      .D       (p2_dl[17]    ),
      .Q       (p3_dl[17]    )
   );
   (* BEL="X2/Y3/lc2" *)
   SB_DFF  dff_2_18 (
      .C       (i_clk         ),
      .D       (p0_dl[19]  ),
      .Q       (p1_dl[18]    )
   );

   (* BEL="X3/Y3/lc2" *)
   SB_DFF  dff_3_18 (
      .C       (i_clk         ),
      .D       (p1_dl[18]    ),
      .Q       (p2_dl[18]    )
   );


   (* BEL="X29/Y3/lc2" *)
   SB_DFF  dff_29_18 (
      .C       (i_clk         ),
      .D       (p2_dl[18]    ),
      .Q       (p3_dl[18]    )
   );
   (* BEL="X2/Y3/lc3" *)
   SB_DFF  dff_2_19 (
      .C       (i_clk         ),
      .D       (p0_dl[20]  ),
      .Q       (p1_dl[19]    )
   );

   (* BEL="X3/Y3/lc3" *)
   SB_DFF  dff_3_19 (
      .C       (i_clk         ),
      .D       (p1_dl[19]    ),
      .Q       (p2_dl[19]    )
   );


   (* BEL="X29/Y3/lc3" *)
   SB_DFF  dff_29_19 (
      .C       (i_clk         ),
      .D       (p2_dl[19]    ),
      .Q       (p3_dl[19]    )
   );
   (* BEL="X2/Y3/lc4" *)
   SB_DFF  dff_2_20 (
      .C       (i_clk         ),
      .D       (p0_dl[21]  ),
      .Q       (p1_dl[20]    )
   );

   (* BEL="X3/Y3/lc4" *)
   SB_DFF  dff_3_20 (
      .C       (i_clk         ),
      .D       (p1_dl[20]    ),
      .Q       (p2_dl[20]    )
   );


   (* BEL="X29/Y3/lc4" *)
   SB_DFF  dff_29_20 (
      .C       (i_clk         ),
      .D       (p2_dl[20]    ),
      .Q       (p3_dl[20]    )
   );
   (* BEL="X2/Y3/lc5" *)
   SB_DFF  dff_2_21 (
      .C       (i_clk         ),
      .D       (p0_dl[22]  ),
      .Q       (p1_dl[21]    )
   );

   (* BEL="X3/Y3/lc5" *)
   SB_DFF  dff_3_21 (
      .C       (i_clk         ),
      .D       (p1_dl[21]    ),
      .Q       (p2_dl[21]    )
   );


   (* BEL="X29/Y3/lc5" *)
   SB_DFF  dff_29_21 (
      .C       (i_clk         ),
      .D       (p2_dl[21]    ),
      .Q       (p3_dl[21]    )
   );
   (* BEL="X2/Y3/lc6" *)
   SB_DFF  dff_2_22 (
      .C       (i_clk         ),
      .D       (p0_dl[23]  ),
      .Q       (p1_dl[22]    )
   );

   (* BEL="X3/Y3/lc6" *)
   SB_DFF  dff_3_22 (
      .C       (i_clk         ),
      .D       (p1_dl[22]    ),
      .Q       (p2_dl[22]    )
   );


   (* BEL="X29/Y3/lc6" *)
   SB_DFF  dff_29_22 (
      .C       (i_clk         ),
      .D       (p2_dl[22]    ),
      .Q       (p3_dl[22]    )
   );
   (* BEL="X2/Y3/lc7" *)
   SB_DFF  dff_2_23 (
      .C       (i_clk         ),
      .D       (p0_dl[24]  ),
      .Q       (p1_dl[23]    )
   );

   (* BEL="X3/Y3/lc7" *)
   SB_DFF  dff_3_23 (
      .C       (i_clk         ),
      .D       (p1_dl[23]    ),
      .Q       (p2_dl[23]    )
   );


   (* BEL="X29/Y3/lc7" *)
   SB_DFF  dff_29_23 (
      .C       (i_clk         ),
      .D       (p2_dl[23]    ),
      .Q       (p3_dl[23]    )
   );
   (* BEL="X2/Y4/lc0" *)
   SB_DFF  dff_2_24 (
      .C       (i_clk         ),
      .D       (p0_dl[25]  ),
      .Q       (p1_dl[24]    )
   );

   (* BEL="X3/Y4/lc0" *)
   SB_DFF  dff_3_24 (
      .C       (i_clk         ),
      .D       (p1_dl[24]    ),
      .Q       (p2_dl[24]    )
   );


   (* BEL="X29/Y4/lc0" *)
   SB_DFF  dff_29_24 (
      .C       (i_clk         ),
      .D       (p2_dl[24]    ),
      .Q       (p3_dl[24]    )
   );
   (* BEL="X2/Y4/lc1" *)
   SB_DFF  dff_2_25 (
      .C       (i_clk         ),
      .D       (p0_dl[26]  ),
      .Q       (p1_dl[25]    )
   );

   (* BEL="X3/Y4/lc1" *)
   SB_DFF  dff_3_25 (
      .C       (i_clk         ),
      .D       (p1_dl[25]    ),
      .Q       (p2_dl[25]    )
   );


   (* BEL="X29/Y4/lc1" *)
   SB_DFF  dff_29_25 (
      .C       (i_clk         ),
      .D       (p2_dl[25]    ),
      .Q       (p3_dl[25]    )
   );
   (* BEL="X2/Y4/lc2" *)
   SB_DFF  dff_2_26 (
      .C       (i_clk         ),
      .D       (p0_dl[27]  ),
      .Q       (p1_dl[26]    )
   );

   (* BEL="X3/Y4/lc2" *)
   SB_DFF  dff_3_26 (
      .C       (i_clk         ),
      .D       (p1_dl[26]    ),
      .Q       (p2_dl[26]    )
   );


   (* BEL="X29/Y4/lc2" *)
   SB_DFF  dff_29_26 (
      .C       (i_clk         ),
      .D       (p2_dl[26]    ),
      .Q       (p3_dl[26]    )
   );
   (* BEL="X2/Y4/lc3" *)
   SB_DFF  dff_2_27 (
      .C       (i_clk         ),
      .D       (p0_dl[28]  ),
      .Q       (p1_dl[27]    )
   );

   (* BEL="X3/Y4/lc3" *)
   SB_DFF  dff_3_27 (
      .C       (i_clk         ),
      .D       (p1_dl[27]    ),
      .Q       (p2_dl[27]    )
   );


   (* BEL="X29/Y4/lc3" *)
   SB_DFF  dff_29_27 (
      .C       (i_clk         ),
      .D       (p2_dl[27]    ),
      .Q       (p3_dl[27]    )
   );
   (* BEL="X2/Y4/lc4" *)
   SB_DFF  dff_2_28 (
      .C       (i_clk         ),
      .D       (p0_dl[29]  ),
      .Q       (p1_dl[28]    )
   );

   (* BEL="X3/Y4/lc4" *)
   SB_DFF  dff_3_28 (
      .C       (i_clk         ),
      .D       (p1_dl[28]    ),
      .Q       (p2_dl[28]    )
   );


   (* BEL="X29/Y4/lc4" *)
   SB_DFF  dff_29_28 (
      .C       (i_clk         ),
      .D       (p2_dl[28]    ),
      .Q       (p3_dl[28]    )
   );
   (* BEL="X2/Y4/lc5" *)
   SB_DFF  dff_2_29 (
      .C       (i_clk         ),
      .D       (p0_dl[30]  ),
      .Q       (p1_dl[29]    )
   );

   (* BEL="X3/Y4/lc5" *)
   SB_DFF  dff_3_29 (
      .C       (i_clk         ),
      .D       (p1_dl[29]    ),
      .Q       (p2_dl[29]    )
   );


   (* BEL="X29/Y4/lc5" *)
   SB_DFF  dff_29_29 (
      .C       (i_clk         ),
      .D       (p2_dl[29]    ),
      .Q       (p3_dl[29]    )
   );
   (* BEL="X2/Y4/lc6" *)
   SB_DFF  dff_2_30 (
      .C       (i_clk         ),
      .D       (p0_dl[31]  ),
      .Q       (p1_dl[30]    )
   );

   (* BEL="X3/Y4/lc6" *)
   SB_DFF  dff_3_30 (
      .C       (i_clk         ),
      .D       (p1_dl[30]    ),
      .Q       (p2_dl[30]    )
   );


   (* BEL="X29/Y4/lc6" *)
   SB_DFF  dff_29_30 (
      .C       (i_clk         ),
      .D       (p2_dl[30]    ),
      .Q       (p3_dl[30]    )
   );
   (* BEL="X2/Y4/lc7" *)
   SB_DFF  dff_2_31 (
      .C       (i_clk         ),
      .D       (p0_dl[32]  ),
      .Q       (p1_dl[31]    )
   );

   (* BEL="X3/Y4/lc7" *)
   SB_DFF  dff_3_31 (
      .C       (i_clk         ),
      .D       (p1_dl[31]    ),
      .Q       (p2_dl[31]    )
   );


   (* BEL="X29/Y4/lc7" *)
   SB_DFF  dff_29_31 (
      .C       (i_clk         ),
      .D       (p2_dl[31]    ),
      .Q       (p3_dl[31]    )
   );
   (* BEL="X2/Y5/lc0" *)
   SB_DFF  dff_2_32 (
      .C       (i_clk         ),
      .D       (p0_dl[33]  ),
      .Q       (p1_dl[32]    )
   );

   (* BEL="X3/Y5/lc0" *)
   SB_DFF  dff_3_32 (
      .C       (i_clk         ),
      .D       (p1_dl[32]    ),
      .Q       (p2_dl[32]    )
   );


   (* BEL="X29/Y5/lc0" *)
   SB_DFF  dff_29_32 (
      .C       (i_clk         ),
      .D       (p2_dl[32]    ),
      .Q       (p3_dl[32]    )
   );
   (* BEL="X2/Y5/lc1" *)
   SB_DFF  dff_2_33 (
      .C       (i_clk         ),
      .D       (p0_dl[34]  ),
      .Q       (p1_dl[33]    )
   );

   (* BEL="X3/Y5/lc1" *)
   SB_DFF  dff_3_33 (
      .C       (i_clk         ),
      .D       (p1_dl[33]    ),
      .Q       (p2_dl[33]    )
   );


   (* BEL="X29/Y5/lc1" *)
   SB_DFF  dff_29_33 (
      .C       (i_clk         ),
      .D       (p2_dl[33]    ),
      .Q       (p3_dl[33]    )
   );
   (* BEL="X2/Y5/lc2" *)
   SB_DFF  dff_2_34 (
      .C       (i_clk         ),
      .D       (p0_dl[35]  ),
      .Q       (p1_dl[34]    )
   );

   (* BEL="X3/Y5/lc2" *)
   SB_DFF  dff_3_34 (
      .C       (i_clk         ),
      .D       (p1_dl[34]    ),
      .Q       (p2_dl[34]    )
   );


   (* BEL="X29/Y5/lc2" *)
   SB_DFF  dff_29_34 (
      .C       (i_clk         ),
      .D       (p2_dl[34]    ),
      .Q       (p3_dl[34]    )
   );
   (* BEL="X2/Y5/lc3" *)
   SB_DFF  dff_2_35 (
      .C       (i_clk         ),
      .D       (p0_dl[36]  ),
      .Q       (p1_dl[35]    )
   );

   (* BEL="X3/Y5/lc3" *)
   SB_DFF  dff_3_35 (
      .C       (i_clk         ),
      .D       (p1_dl[35]    ),
      .Q       (p2_dl[35]    )
   );


   (* BEL="X29/Y5/lc3" *)
   SB_DFF  dff_29_35 (
      .C       (i_clk         ),
      .D       (p2_dl[35]    ),
      .Q       (p3_dl[35]    )
   );
   (* BEL="X2/Y5/lc4" *)
   SB_DFF  dff_2_36 (
      .C       (i_clk         ),
      .D       (p0_dl[37]  ),
      .Q       (p1_dl[36]    )
   );

   (* BEL="X3/Y5/lc4" *)
   SB_DFF  dff_3_36 (
      .C       (i_clk         ),
      .D       (p1_dl[36]    ),
      .Q       (p2_dl[36]    )
   );


   (* BEL="X29/Y5/lc4" *)
   SB_DFF  dff_29_36 (
      .C       (i_clk         ),
      .D       (p2_dl[36]    ),
      .Q       (p3_dl[36]    )
   );
   (* BEL="X2/Y5/lc5" *)
   SB_DFF  dff_2_37 (
      .C       (i_clk         ),
      .D       (p0_dl[38]  ),
      .Q       (p1_dl[37]    )
   );

   (* BEL="X3/Y5/lc5" *)
   SB_DFF  dff_3_37 (
      .C       (i_clk         ),
      .D       (p1_dl[37]    ),
      .Q       (p2_dl[37]    )
   );


   (* BEL="X29/Y5/lc5" *)
   SB_DFF  dff_29_37 (
      .C       (i_clk         ),
      .D       (p2_dl[37]    ),
      .Q       (p3_dl[37]    )
   );
   (* BEL="X2/Y5/lc6" *)
   SB_DFF  dff_2_38 (
      .C       (i_clk         ),
      .D       (p0_dl[39]  ),
      .Q       (p1_dl[38]    )
   );

   (* BEL="X3/Y5/lc6" *)
   SB_DFF  dff_3_38 (
      .C       (i_clk         ),
      .D       (p1_dl[38]    ),
      .Q       (p2_dl[38]    )
   );


   (* BEL="X29/Y5/lc6" *)
   SB_DFF  dff_29_38 (
      .C       (i_clk         ),
      .D       (p2_dl[38]    ),
      .Q       (p3_dl[38]    )
   );
   (* BEL="X2/Y5/lc7" *)
   SB_DFF  dff_2_39 (
      .C       (i_clk         ),
      .D       (p0_dl[40]  ),
      .Q       (p1_dl[39]    )
   );

   (* BEL="X3/Y5/lc7" *)
   SB_DFF  dff_3_39 (
      .C       (i_clk         ),
      .D       (p1_dl[39]    ),
      .Q       (p2_dl[39]    )
   );


   (* BEL="X29/Y5/lc7" *)
   SB_DFF  dff_29_39 (
      .C       (i_clk         ),
      .D       (p2_dl[39]    ),
      .Q       (p3_dl[39]    )
   );
   (* BEL="X2/Y6/lc0" *)
   SB_DFF  dff_2_40 (
      .C       (i_clk         ),
      .D       (p0_dl[41]  ),
      .Q       (p1_dl[40]    )
   );

   (* BEL="X3/Y6/lc0" *)
   SB_DFF  dff_3_40 (
      .C       (i_clk         ),
      .D       (p1_dl[40]    ),
      .Q       (p2_dl[40]    )
   );


   (* BEL="X29/Y6/lc0" *)
   SB_DFF  dff_29_40 (
      .C       (i_clk         ),
      .D       (p2_dl[40]    ),
      .Q       (p3_dl[40]    )
   );
   (* BEL="X2/Y6/lc1" *)
   SB_DFF  dff_2_41 (
      .C       (i_clk         ),
      .D       (p0_dl[42]  ),
      .Q       (p1_dl[41]    )
   );

   (* BEL="X3/Y6/lc1" *)
   SB_DFF  dff_3_41 (
      .C       (i_clk         ),
      .D       (p1_dl[41]    ),
      .Q       (p2_dl[41]    )
   );


   (* BEL="X29/Y6/lc1" *)
   SB_DFF  dff_29_41 (
      .C       (i_clk         ),
      .D       (p2_dl[41]    ),
      .Q       (p3_dl[41]    )
   );
   (* BEL="X2/Y6/lc2" *)
   SB_DFF  dff_2_42 (
      .C       (i_clk         ),
      .D       (p0_dl[43]  ),
      .Q       (p1_dl[42]    )
   );

   (* BEL="X3/Y6/lc2" *)
   SB_DFF  dff_3_42 (
      .C       (i_clk         ),
      .D       (p1_dl[42]    ),
      .Q       (p2_dl[42]    )
   );


   (* BEL="X29/Y6/lc2" *)
   SB_DFF  dff_29_42 (
      .C       (i_clk         ),
      .D       (p2_dl[42]    ),
      .Q       (p3_dl[42]    )
   );
   (* BEL="X2/Y6/lc3" *)
   SB_DFF  dff_2_43 (
      .C       (i_clk         ),
      .D       (p0_dl[44]  ),
      .Q       (p1_dl[43]    )
   );

   (* BEL="X3/Y6/lc3" *)
   SB_DFF  dff_3_43 (
      .C       (i_clk         ),
      .D       (p1_dl[43]    ),
      .Q       (p2_dl[43]    )
   );


   (* BEL="X29/Y6/lc3" *)
   SB_DFF  dff_29_43 (
      .C       (i_clk         ),
      .D       (p2_dl[43]    ),
      .Q       (p3_dl[43]    )
   );
   (* BEL="X2/Y6/lc4" *)
   SB_DFF  dff_2_44 (
      .C       (i_clk         ),
      .D       (p0_dl[45]  ),
      .Q       (p1_dl[44]    )
   );

   (* BEL="X3/Y6/lc4" *)
   SB_DFF  dff_3_44 (
      .C       (i_clk         ),
      .D       (p1_dl[44]    ),
      .Q       (p2_dl[44]    )
   );


   (* BEL="X29/Y6/lc4" *)
   SB_DFF  dff_29_44 (
      .C       (i_clk         ),
      .D       (p2_dl[44]    ),
      .Q       (p3_dl[44]    )
   );
   (* BEL="X2/Y6/lc5" *)
   SB_DFF  dff_2_45 (
      .C       (i_clk         ),
      .D       (p0_dl[46]  ),
      .Q       (p1_dl[45]    )
   );

   (* BEL="X3/Y6/lc5" *)
   SB_DFF  dff_3_45 (
      .C       (i_clk         ),
      .D       (p1_dl[45]    ),
      .Q       (p2_dl[45]    )
   );


   (* BEL="X29/Y6/lc5" *)
   SB_DFF  dff_29_45 (
      .C       (i_clk         ),
      .D       (p2_dl[45]    ),
      .Q       (p3_dl[45]    )
   );
   (* BEL="X2/Y6/lc6" *)
   SB_DFF  dff_2_46 (
      .C       (i_clk         ),
      .D       (p0_dl[47]  ),
      .Q       (p1_dl[46]    )
   );

   (* BEL="X3/Y6/lc6" *)
   SB_DFF  dff_3_46 (
      .C       (i_clk         ),
      .D       (p1_dl[46]    ),
      .Q       (p2_dl[46]    )
   );


   (* BEL="X29/Y6/lc6" *)
   SB_DFF  dff_29_46 (
      .C       (i_clk         ),
      .D       (p2_dl[46]    ),
      .Q       (p3_dl[46]    )
   );
   (* BEL="X2/Y6/lc7" *)
   SB_DFF  dff_2_47 (
      .C       (i_clk         ),
      .D       (p0_dl[48]  ),
      .Q       (p1_dl[47]    )
   );

   (* BEL="X3/Y6/lc7" *)
   SB_DFF  dff_3_47 (
      .C       (i_clk         ),
      .D       (p1_dl[47]    ),
      .Q       (p2_dl[47]    )
   );


   (* BEL="X29/Y6/lc7" *)
   SB_DFF  dff_29_47 (
      .C       (i_clk         ),
      .D       (p2_dl[47]    ),
      .Q       (p3_dl[47]    )
   );
   (* BEL="X2/Y7/lc0" *)
   SB_DFF  dff_2_48 (
      .C       (i_clk         ),
      .D       (p0_dl[49]  ),
      .Q       (p1_dl[48]    )
   );

   (* BEL="X3/Y7/lc0" *)
   SB_DFF  dff_3_48 (
      .C       (i_clk         ),
      .D       (p1_dl[48]    ),
      .Q       (p2_dl[48]    )
   );


   (* BEL="X29/Y7/lc0" *)
   SB_DFF  dff_29_48 (
      .C       (i_clk         ),
      .D       (p2_dl[48]    ),
      .Q       (p3_dl[48]    )
   );
   (* BEL="X2/Y7/lc1" *)
   SB_DFF  dff_2_49 (
      .C       (i_clk         ),
      .D       (p0_dl[50]  ),
      .Q       (p1_dl[49]    )
   );

   (* BEL="X3/Y7/lc1" *)
   SB_DFF  dff_3_49 (
      .C       (i_clk         ),
      .D       (p1_dl[49]    ),
      .Q       (p2_dl[49]    )
   );


   (* BEL="X29/Y7/lc1" *)
   SB_DFF  dff_29_49 (
      .C       (i_clk         ),
      .D       (p2_dl[49]    ),
      .Q       (p3_dl[49]    )
   );
   (* BEL="X2/Y7/lc2" *)
   SB_DFF  dff_2_50 (
      .C       (i_clk         ),
      .D       (p0_dl[51]  ),
      .Q       (p1_dl[50]    )
   );

   (* BEL="X3/Y7/lc2" *)
   SB_DFF  dff_3_50 (
      .C       (i_clk         ),
      .D       (p1_dl[50]    ),
      .Q       (p2_dl[50]    )
   );


   (* BEL="X29/Y7/lc2" *)
   SB_DFF  dff_29_50 (
      .C       (i_clk         ),
      .D       (p2_dl[50]    ),
      .Q       (p3_dl[50]    )
   );
   (* BEL="X2/Y7/lc3" *)
   SB_DFF  dff_2_51 (
      .C       (i_clk         ),
      .D       (p0_dl[52]  ),
      .Q       (p1_dl[51]    )
   );

   (* BEL="X3/Y7/lc3" *)
   SB_DFF  dff_3_51 (
      .C       (i_clk         ),
      .D       (p1_dl[51]    ),
      .Q       (p2_dl[51]    )
   );


   (* BEL="X29/Y7/lc3" *)
   SB_DFF  dff_29_51 (
      .C       (i_clk         ),
      .D       (p2_dl[51]    ),
      .Q       (p3_dl[51]    )
   );
   (* BEL="X2/Y7/lc4" *)
   SB_DFF  dff_2_52 (
      .C       (i_clk         ),
      .D       (p0_dl[53]  ),
      .Q       (p1_dl[52]    )
   );

   (* BEL="X3/Y7/lc4" *)
   SB_DFF  dff_3_52 (
      .C       (i_clk         ),
      .D       (p1_dl[52]    ),
      .Q       (p2_dl[52]    )
   );


   (* BEL="X29/Y7/lc4" *)
   SB_DFF  dff_29_52 (
      .C       (i_clk         ),
      .D       (p2_dl[52]    ),
      .Q       (p3_dl[52]    )
   );
   (* BEL="X2/Y7/lc5" *)
   SB_DFF  dff_2_53 (
      .C       (i_clk         ),
      .D       (p0_dl[54]  ),
      .Q       (p1_dl[53]    )
   );

   (* BEL="X3/Y7/lc5" *)
   SB_DFF  dff_3_53 (
      .C       (i_clk         ),
      .D       (p1_dl[53]    ),
      .Q       (p2_dl[53]    )
   );


   (* BEL="X29/Y7/lc5" *)
   SB_DFF  dff_29_53 (
      .C       (i_clk         ),
      .D       (p2_dl[53]    ),
      .Q       (p3_dl[53]    )
   );
   (* BEL="X2/Y7/lc6" *)
   SB_DFF  dff_2_54 (
      .C       (i_clk         ),
      .D       (p0_dl[55]  ),
      .Q       (p1_dl[54]    )
   );

   (* BEL="X3/Y7/lc6" *)
   SB_DFF  dff_3_54 (
      .C       (i_clk         ),
      .D       (p1_dl[54]    ),
      .Q       (p2_dl[54]    )
   );


   (* BEL="X29/Y7/lc6" *)
   SB_DFF  dff_29_54 (
      .C       (i_clk         ),
      .D       (p2_dl[54]    ),
      .Q       (p3_dl[54]    )
   );
   (* BEL="X2/Y7/lc7" *)
   SB_DFF  dff_2_55 (
      .C       (i_clk         ),
      .D       (p0_dl[56]  ),
      .Q       (p1_dl[55]    )
   );

   (* BEL="X3/Y7/lc7" *)
   SB_DFF  dff_3_55 (
      .C       (i_clk         ),
      .D       (p1_dl[55]    ),
      .Q       (p2_dl[55]    )
   );


   (* BEL="X29/Y7/lc7" *)
   SB_DFF  dff_29_55 (
      .C       (i_clk         ),
      .D       (p2_dl[55]    ),
      .Q       (p3_dl[55]    )
   );
   (* BEL="X2/Y8/lc0" *)
   SB_DFF  dff_2_56 (
      .C       (i_clk         ),
      .D       (p0_dl[57]  ),
      .Q       (p1_dl[56]    )
   );

   (* BEL="X3/Y8/lc0" *)
   SB_DFF  dff_3_56 (
      .C       (i_clk         ),
      .D       (p1_dl[56]    ),
      .Q       (p2_dl[56]    )
   );


   (* BEL="X29/Y8/lc0" *)
   SB_DFF  dff_29_56 (
      .C       (i_clk         ),
      .D       (p2_dl[56]    ),
      .Q       (p3_dl[56]    )
   );
   (* BEL="X2/Y8/lc1" *)
   SB_DFF  dff_2_57 (
      .C       (i_clk         ),
      .D       (p0_dl[58]  ),
      .Q       (p1_dl[57]    )
   );

   (* BEL="X3/Y8/lc1" *)
   SB_DFF  dff_3_57 (
      .C       (i_clk         ),
      .D       (p1_dl[57]    ),
      .Q       (p2_dl[57]    )
   );


   (* BEL="X29/Y8/lc1" *)
   SB_DFF  dff_29_57 (
      .C       (i_clk         ),
      .D       (p2_dl[57]    ),
      .Q       (p3_dl[57]    )
   );
   (* BEL="X2/Y8/lc2" *)
   SB_DFF  dff_2_58 (
      .C       (i_clk         ),
      .D       (p0_dl[59]  ),
      .Q       (p1_dl[58]    )
   );

   (* BEL="X3/Y8/lc2" *)
   SB_DFF  dff_3_58 (
      .C       (i_clk         ),
      .D       (p1_dl[58]    ),
      .Q       (p2_dl[58]    )
   );


   (* BEL="X29/Y8/lc2" *)
   SB_DFF  dff_29_58 (
      .C       (i_clk         ),
      .D       (p2_dl[58]    ),
      .Q       (p3_dl[58]    )
   );
   (* BEL="X2/Y8/lc3" *)
   SB_DFF  dff_2_59 (
      .C       (i_clk         ),
      .D       (p0_dl[60]  ),
      .Q       (p1_dl[59]    )
   );

   (* BEL="X3/Y8/lc3" *)
   SB_DFF  dff_3_59 (
      .C       (i_clk         ),
      .D       (p1_dl[59]    ),
      .Q       (p2_dl[59]    )
   );


   (* BEL="X29/Y8/lc3" *)
   SB_DFF  dff_29_59 (
      .C       (i_clk         ),
      .D       (p2_dl[59]    ),
      .Q       (p3_dl[59]    )
   );
   (* BEL="X2/Y8/lc4" *)
   SB_DFF  dff_2_60 (
      .C       (i_clk         ),
      .D       (p0_dl[61]  ),
      .Q       (p1_dl[60]    )
   );

   (* BEL="X3/Y8/lc4" *)
   SB_DFF  dff_3_60 (
      .C       (i_clk         ),
      .D       (p1_dl[60]    ),
      .Q       (p2_dl[60]    )
   );


   (* BEL="X29/Y8/lc4" *)
   SB_DFF  dff_29_60 (
      .C       (i_clk         ),
      .D       (p2_dl[60]    ),
      .Q       (p3_dl[60]    )
   );
   (* BEL="X2/Y8/lc5" *)
   SB_DFF  dff_2_61 (
      .C       (i_clk         ),
      .D       (p0_dl[62]  ),
      .Q       (p1_dl[61]    )
   );

   (* BEL="X3/Y8/lc5" *)
   SB_DFF  dff_3_61 (
      .C       (i_clk         ),
      .D       (p1_dl[61]    ),
      .Q       (p2_dl[61]    )
   );


   (* BEL="X29/Y8/lc5" *)
   SB_DFF  dff_29_61 (
      .C       (i_clk         ),
      .D       (p2_dl[61]    ),
      .Q       (p3_dl[61]    )
   );
   (* BEL="X2/Y8/lc6" *)
   SB_DFF  dff_2_62 (
      .C       (i_clk         ),
      .D       (p0_dl[63]  ),
      .Q       (p1_dl[62]    )
   );

   (* BEL="X3/Y8/lc6" *)
   SB_DFF  dff_3_62 (
      .C       (i_clk         ),
      .D       (p1_dl[62]    ),
      .Q       (p2_dl[62]    )
   );


   (* BEL="X29/Y8/lc6" *)
   SB_DFF  dff_29_62 (
      .C       (i_clk         ),
      .D       (p2_dl[62]    ),
      .Q       (p3_dl[62]    )
   );
   (* BEL="X2/Y8/lc7" *)
   SB_DFF  dff_2_63 (
      .C       (i_clk         ),
      .D       (p0_dl[64]  ),
      .Q       (p1_dl[63]    )
   );

   (* BEL="X3/Y8/lc7" *)
   SB_DFF  dff_3_63 (
      .C       (i_clk         ),
      .D       (p1_dl[63]    ),
      .Q       (p2_dl[63]    )
   );


   (* BEL="X29/Y8/lc7" *)
   SB_DFF  dff_29_63 (
      .C       (i_clk         ),
      .D       (p2_dl[63]    ),
      .Q       (p3_dl[63]    )
   );
   (* BEL="X2/Y9/lc0" *)
   SB_DFF  dff_2_64 (
      .C       (i_clk         ),
      .D       (p0_dl[65]  ),
      .Q       (p1_dl[64]    )
   );

   (* BEL="X3/Y9/lc0" *)
   SB_DFF  dff_3_64 (
      .C       (i_clk         ),
      .D       (p1_dl[64]    ),
      .Q       (p2_dl[64]    )
   );


   (* BEL="X29/Y9/lc0" *)
   SB_DFF  dff_29_64 (
      .C       (i_clk         ),
      .D       (p2_dl[64]    ),
      .Q       (p3_dl[64]    )
   );
   (* BEL="X2/Y9/lc1" *)
   SB_DFF  dff_2_65 (
      .C       (i_clk         ),
      .D       (p0_dl[66]  ),
      .Q       (p1_dl[65]    )
   );

   (* BEL="X3/Y9/lc1" *)
   SB_DFF  dff_3_65 (
      .C       (i_clk         ),
      .D       (p1_dl[65]    ),
      .Q       (p2_dl[65]    )
   );


   (* BEL="X29/Y9/lc1" *)
   SB_DFF  dff_29_65 (
      .C       (i_clk         ),
      .D       (p2_dl[65]    ),
      .Q       (p3_dl[65]    )
   );
   (* BEL="X2/Y9/lc2" *)
   SB_DFF  dff_2_66 (
      .C       (i_clk         ),
      .D       (p0_dl[67]  ),
      .Q       (p1_dl[66]    )
   );

   (* BEL="X3/Y9/lc2" *)
   SB_DFF  dff_3_66 (
      .C       (i_clk         ),
      .D       (p1_dl[66]    ),
      .Q       (p2_dl[66]    )
   );


   (* BEL="X29/Y9/lc2" *)
   SB_DFF  dff_29_66 (
      .C       (i_clk         ),
      .D       (p2_dl[66]    ),
      .Q       (p3_dl[66]    )
   );
   (* BEL="X2/Y9/lc3" *)
   SB_DFF  dff_2_67 (
      .C       (i_clk         ),
      .D       (p0_dl[68]  ),
      .Q       (p1_dl[67]    )
   );

   (* BEL="X3/Y9/lc3" *)
   SB_DFF  dff_3_67 (
      .C       (i_clk         ),
      .D       (p1_dl[67]    ),
      .Q       (p2_dl[67]    )
   );


   (* BEL="X29/Y9/lc3" *)
   SB_DFF  dff_29_67 (
      .C       (i_clk         ),
      .D       (p2_dl[67]    ),
      .Q       (p3_dl[67]    )
   );
   (* BEL="X2/Y9/lc4" *)
   SB_DFF  dff_2_68 (
      .C       (i_clk         ),
      .D       (p0_dl[69]  ),
      .Q       (p1_dl[68]    )
   );

   (* BEL="X3/Y9/lc4" *)
   SB_DFF  dff_3_68 (
      .C       (i_clk         ),
      .D       (p1_dl[68]    ),
      .Q       (p2_dl[68]    )
   );


   (* BEL="X29/Y9/lc4" *)
   SB_DFF  dff_29_68 (
      .C       (i_clk         ),
      .D       (p2_dl[68]    ),
      .Q       (p3_dl[68]    )
   );
   (* BEL="X2/Y9/lc5" *)
   SB_DFF  dff_2_69 (
      .C       (i_clk         ),
      .D       (p0_dl[70]  ),
      .Q       (p1_dl[69]    )
   );

   (* BEL="X3/Y9/lc5" *)
   SB_DFF  dff_3_69 (
      .C       (i_clk         ),
      .D       (p1_dl[69]    ),
      .Q       (p2_dl[69]    )
   );


   (* BEL="X29/Y9/lc5" *)
   SB_DFF  dff_29_69 (
      .C       (i_clk         ),
      .D       (p2_dl[69]    ),
      .Q       (p3_dl[69]    )
   );
   (* BEL="X2/Y9/lc6" *)
   SB_DFF  dff_2_70 (
      .C       (i_clk         ),
      .D       (p0_dl[71]  ),
      .Q       (p1_dl[70]    )
   );

   (* BEL="X3/Y9/lc6" *)
   SB_DFF  dff_3_70 (
      .C       (i_clk         ),
      .D       (p1_dl[70]    ),
      .Q       (p2_dl[70]    )
   );


   (* BEL="X29/Y9/lc6" *)
   SB_DFF  dff_29_70 (
      .C       (i_clk         ),
      .D       (p2_dl[70]    ),
      .Q       (p3_dl[70]    )
   );
   (* BEL="X2/Y9/lc7" *)
   SB_DFF  dff_2_71 (
      .C       (i_clk         ),
      .D       (p0_dl[72]  ),
      .Q       (p1_dl[71]    )
   );

   (* BEL="X3/Y9/lc7" *)
   SB_DFF  dff_3_71 (
      .C       (i_clk         ),
      .D       (p1_dl[71]    ),
      .Q       (p2_dl[71]    )
   );


   (* BEL="X29/Y9/lc7" *)
   SB_DFF  dff_29_71 (
      .C       (i_clk         ),
      .D       (p2_dl[71]    ),
      .Q       (p3_dl[71]    )
   );
   (* BEL="X2/Y10/lc0" *)
   SB_DFF  dff_2_72 (
      .C       (i_clk         ),
      .D       (p0_dl[73]  ),
      .Q       (p1_dl[72]    )
   );

   (* BEL="X3/Y10/lc0" *)
   SB_DFF  dff_3_72 (
      .C       (i_clk         ),
      .D       (p1_dl[72]    ),
      .Q       (p2_dl[72]    )
   );


   (* BEL="X29/Y10/lc0" *)
   SB_DFF  dff_29_72 (
      .C       (i_clk         ),
      .D       (p2_dl[72]    ),
      .Q       (p3_dl[72]    )
   );
   (* BEL="X2/Y10/lc1" *)
   SB_DFF  dff_2_73 (
      .C       (i_clk         ),
      .D       (p0_dl[74]  ),
      .Q       (p1_dl[73]    )
   );

   (* BEL="X3/Y10/lc1" *)
   SB_DFF  dff_3_73 (
      .C       (i_clk         ),
      .D       (p1_dl[73]    ),
      .Q       (p2_dl[73]    )
   );


   (* BEL="X29/Y10/lc1" *)
   SB_DFF  dff_29_73 (
      .C       (i_clk         ),
      .D       (p2_dl[73]    ),
      .Q       (p3_dl[73]    )
   );
   (* BEL="X2/Y10/lc2" *)
   SB_DFF  dff_2_74 (
      .C       (i_clk         ),
      .D       (p0_dl[75]  ),
      .Q       (p1_dl[74]    )
   );

   (* BEL="X3/Y10/lc2" *)
   SB_DFF  dff_3_74 (
      .C       (i_clk         ),
      .D       (p1_dl[74]    ),
      .Q       (p2_dl[74]    )
   );


   (* BEL="X29/Y10/lc2" *)
   SB_DFF  dff_29_74 (
      .C       (i_clk         ),
      .D       (p2_dl[74]    ),
      .Q       (p3_dl[74]    )
   );
   (* BEL="X2/Y10/lc3" *)
   SB_DFF  dff_2_75 (
      .C       (i_clk         ),
      .D       (p0_dl[76]  ),
      .Q       (p1_dl[75]    )
   );

   (* BEL="X3/Y10/lc3" *)
   SB_DFF  dff_3_75 (
      .C       (i_clk         ),
      .D       (p1_dl[75]    ),
      .Q       (p2_dl[75]    )
   );


   (* BEL="X29/Y10/lc3" *)
   SB_DFF  dff_29_75 (
      .C       (i_clk         ),
      .D       (p2_dl[75]    ),
      .Q       (p3_dl[75]    )
   );
   (* BEL="X2/Y10/lc4" *)
   SB_DFF  dff_2_76 (
      .C       (i_clk         ),
      .D       (p0_dl[77]  ),
      .Q       (p1_dl[76]    )
   );

   (* BEL="X3/Y10/lc4" *)
   SB_DFF  dff_3_76 (
      .C       (i_clk         ),
      .D       (p1_dl[76]    ),
      .Q       (p2_dl[76]    )
   );


   (* BEL="X29/Y10/lc4" *)
   SB_DFF  dff_29_76 (
      .C       (i_clk         ),
      .D       (p2_dl[76]    ),
      .Q       (p3_dl[76]    )
   );
   (* BEL="X2/Y10/lc5" *)
   SB_DFF  dff_2_77 (
      .C       (i_clk         ),
      .D       (p0_dl[78]  ),
      .Q       (p1_dl[77]    )
   );

   (* BEL="X3/Y10/lc5" *)
   SB_DFF  dff_3_77 (
      .C       (i_clk         ),
      .D       (p1_dl[77]    ),
      .Q       (p2_dl[77]    )
   );


   (* BEL="X29/Y10/lc5" *)
   SB_DFF  dff_29_77 (
      .C       (i_clk         ),
      .D       (p2_dl[77]    ),
      .Q       (p3_dl[77]    )
   );
   (* BEL="X2/Y10/lc6" *)
   SB_DFF  dff_2_78 (
      .C       (i_clk         ),
      .D       (p0_dl[79]  ),
      .Q       (p1_dl[78]    )
   );

   (* BEL="X3/Y10/lc6" *)
   SB_DFF  dff_3_78 (
      .C       (i_clk         ),
      .D       (p1_dl[78]    ),
      .Q       (p2_dl[78]    )
   );


   (* BEL="X29/Y10/lc6" *)
   SB_DFF  dff_29_78 (
      .C       (i_clk         ),
      .D       (p2_dl[78]    ),
      .Q       (p3_dl[78]    )
   );
   (* BEL="X2/Y10/lc7" *)
   SB_DFF  dff_2_79 (
      .C       (i_clk         ),
      .D       (p0_dl[80]  ),
      .Q       (p1_dl[79]    )
   );

   (* BEL="X3/Y10/lc7" *)
   SB_DFF  dff_3_79 (
      .C       (i_clk         ),
      .D       (p1_dl[79]    ),
      .Q       (p2_dl[79]    )
   );


   (* BEL="X29/Y10/lc7" *)
   SB_DFF  dff_29_79 (
      .C       (i_clk         ),
      .D       (p2_dl[79]    ),
      .Q       (p3_dl[79]    )
   );
   (* BEL="X2/Y11/lc0" *)
   SB_DFF  dff_2_80 (
      .C       (i_clk         ),
      .D       (p0_dl[81]  ),
      .Q       (p1_dl[80]    )
   );

   (* BEL="X3/Y11/lc0" *)
   SB_DFF  dff_3_80 (
      .C       (i_clk         ),
      .D       (p1_dl[80]    ),
      .Q       (p2_dl[80]    )
   );


   (* BEL="X29/Y11/lc0" *)
   SB_DFF  dff_29_80 (
      .C       (i_clk         ),
      .D       (p2_dl[80]    ),
      .Q       (p3_dl[80]    )
   );
   (* BEL="X2/Y11/lc1" *)
   SB_DFF  dff_2_81 (
      .C       (i_clk         ),
      .D       (p0_dl[82]  ),
      .Q       (p1_dl[81]    )
   );

   (* BEL="X3/Y11/lc1" *)
   SB_DFF  dff_3_81 (
      .C       (i_clk         ),
      .D       (p1_dl[81]    ),
      .Q       (p2_dl[81]    )
   );


   (* BEL="X29/Y11/lc1" *)
   SB_DFF  dff_29_81 (
      .C       (i_clk         ),
      .D       (p2_dl[81]    ),
      .Q       (p3_dl[81]    )
   );
   (* BEL="X2/Y11/lc2" *)
   SB_DFF  dff_2_82 (
      .C       (i_clk         ),
      .D       (p0_dl[83]  ),
      .Q       (p1_dl[82]    )
   );

   (* BEL="X3/Y11/lc2" *)
   SB_DFF  dff_3_82 (
      .C       (i_clk         ),
      .D       (p1_dl[82]    ),
      .Q       (p2_dl[82]    )
   );


   (* BEL="X29/Y11/lc2" *)
   SB_DFF  dff_29_82 (
      .C       (i_clk         ),
      .D       (p2_dl[82]    ),
      .Q       (p3_dl[82]    )
   );
   (* BEL="X2/Y11/lc3" *)
   SB_DFF  dff_2_83 (
      .C       (i_clk         ),
      .D       (p0_dl[84]  ),
      .Q       (p1_dl[83]    )
   );

   (* BEL="X3/Y11/lc3" *)
   SB_DFF  dff_3_83 (
      .C       (i_clk         ),
      .D       (p1_dl[83]    ),
      .Q       (p2_dl[83]    )
   );


   (* BEL="X29/Y11/lc3" *)
   SB_DFF  dff_29_83 (
      .C       (i_clk         ),
      .D       (p2_dl[83]    ),
      .Q       (p3_dl[83]    )
   );
   (* BEL="X2/Y11/lc4" *)
   SB_DFF  dff_2_84 (
      .C       (i_clk         ),
      .D       (p0_dl[85]  ),
      .Q       (p1_dl[84]    )
   );

   (* BEL="X3/Y11/lc4" *)
   SB_DFF  dff_3_84 (
      .C       (i_clk         ),
      .D       (p1_dl[84]    ),
      .Q       (p2_dl[84]    )
   );


   (* BEL="X29/Y11/lc4" *)
   SB_DFF  dff_29_84 (
      .C       (i_clk         ),
      .D       (p2_dl[84]    ),
      .Q       (p3_dl[84]    )
   );
   (* BEL="X2/Y11/lc5" *)
   SB_DFF  dff_2_85 (
      .C       (i_clk         ),
      .D       (p0_dl[86]  ),
      .Q       (p1_dl[85]    )
   );

   (* BEL="X3/Y11/lc5" *)
   SB_DFF  dff_3_85 (
      .C       (i_clk         ),
      .D       (p1_dl[85]    ),
      .Q       (p2_dl[85]    )
   );


   (* BEL="X29/Y11/lc5" *)
   SB_DFF  dff_29_85 (
      .C       (i_clk         ),
      .D       (p2_dl[85]    ),
      .Q       (p3_dl[85]    )
   );
   (* BEL="X2/Y11/lc6" *)
   SB_DFF  dff_2_86 (
      .C       (i_clk         ),
      .D       (p0_dl[87]  ),
      .Q       (p1_dl[86]    )
   );

   (* BEL="X3/Y11/lc6" *)
   SB_DFF  dff_3_86 (
      .C       (i_clk         ),
      .D       (p1_dl[86]    ),
      .Q       (p2_dl[86]    )
   );


   (* BEL="X29/Y11/lc6" *)
   SB_DFF  dff_29_86 (
      .C       (i_clk         ),
      .D       (p2_dl[86]    ),
      .Q       (p3_dl[86]    )
   );
   (* BEL="X2/Y11/lc7" *)
   SB_DFF  dff_2_87 (
      .C       (i_clk         ),
      .D       (p0_dl[88]  ),
      .Q       (p1_dl[87]    )
   );

   (* BEL="X3/Y11/lc7" *)
   SB_DFF  dff_3_87 (
      .C       (i_clk         ),
      .D       (p1_dl[87]    ),
      .Q       (p2_dl[87]    )
   );


   (* BEL="X29/Y11/lc7" *)
   SB_DFF  dff_29_87 (
      .C       (i_clk         ),
      .D       (p2_dl[87]    ),
      .Q       (p3_dl[87]    )
   );
   (* BEL="X2/Y12/lc0" *)
   SB_DFF  dff_2_88 (
      .C       (i_clk         ),
      .D       (p0_dl[89]  ),
      .Q       (p1_dl[88]    )
   );

   (* BEL="X3/Y12/lc0" *)
   SB_DFF  dff_3_88 (
      .C       (i_clk         ),
      .D       (p1_dl[88]    ),
      .Q       (p2_dl[88]    )
   );


   (* BEL="X29/Y12/lc0" *)
   SB_DFF  dff_29_88 (
      .C       (i_clk         ),
      .D       (p2_dl[88]    ),
      .Q       (p3_dl[88]    )
   );
   (* BEL="X2/Y12/lc1" *)
   SB_DFF  dff_2_89 (
      .C       (i_clk         ),
      .D       (p0_dl[90]  ),
      .Q       (p1_dl[89]    )
   );

   (* BEL="X3/Y12/lc1" *)
   SB_DFF  dff_3_89 (
      .C       (i_clk         ),
      .D       (p1_dl[89]    ),
      .Q       (p2_dl[89]    )
   );


   (* BEL="X29/Y12/lc1" *)
   SB_DFF  dff_29_89 (
      .C       (i_clk         ),
      .D       (p2_dl[89]    ),
      .Q       (p3_dl[89]    )
   );
   (* BEL="X2/Y12/lc2" *)
   SB_DFF  dff_2_90 (
      .C       (i_clk         ),
      .D       (p0_dl[91]  ),
      .Q       (p1_dl[90]    )
   );

   (* BEL="X3/Y12/lc2" *)
   SB_DFF  dff_3_90 (
      .C       (i_clk         ),
      .D       (p1_dl[90]    ),
      .Q       (p2_dl[90]    )
   );


   (* BEL="X29/Y12/lc2" *)
   SB_DFF  dff_29_90 (
      .C       (i_clk         ),
      .D       (p2_dl[90]    ),
      .Q       (p3_dl[90]    )
   );
   (* BEL="X2/Y12/lc3" *)
   SB_DFF  dff_2_91 (
      .C       (i_clk         ),
      .D       (p0_dl[92]  ),
      .Q       (p1_dl[91]    )
   );

   (* BEL="X3/Y12/lc3" *)
   SB_DFF  dff_3_91 (
      .C       (i_clk         ),
      .D       (p1_dl[91]    ),
      .Q       (p2_dl[91]    )
   );


   (* BEL="X29/Y12/lc3" *)
   SB_DFF  dff_29_91 (
      .C       (i_clk         ),
      .D       (p2_dl[91]    ),
      .Q       (p3_dl[91]    )
   );
   (* BEL="X2/Y12/lc4" *)
   SB_DFF  dff_2_92 (
      .C       (i_clk         ),
      .D       (p0_dl[93]  ),
      .Q       (p1_dl[92]    )
   );

   (* BEL="X3/Y12/lc4" *)
   SB_DFF  dff_3_92 (
      .C       (i_clk         ),
      .D       (p1_dl[92]    ),
      .Q       (p2_dl[92]    )
   );


   (* BEL="X29/Y12/lc4" *)
   SB_DFF  dff_29_92 (
      .C       (i_clk         ),
      .D       (p2_dl[92]    ),
      .Q       (p3_dl[92]    )
   );
   (* BEL="X2/Y12/lc5" *)
   SB_DFF  dff_2_93 (
      .C       (i_clk         ),
      .D       (p0_dl[94]  ),
      .Q       (p1_dl[93]    )
   );

   (* BEL="X3/Y12/lc5" *)
   SB_DFF  dff_3_93 (
      .C       (i_clk         ),
      .D       (p1_dl[93]    ),
      .Q       (p2_dl[93]    )
   );


   (* BEL="X29/Y12/lc5" *)
   SB_DFF  dff_29_93 (
      .C       (i_clk         ),
      .D       (p2_dl[93]    ),
      .Q       (p3_dl[93]    )
   );
   (* BEL="X2/Y12/lc6" *)
   SB_DFF  dff_2_94 (
      .C       (i_clk         ),
      .D       (p0_dl[95]  ),
      .Q       (p1_dl[94]    )
   );

   (* BEL="X3/Y12/lc6" *)
   SB_DFF  dff_3_94 (
      .C       (i_clk         ),
      .D       (p1_dl[94]    ),
      .Q       (p2_dl[94]    )
   );


   (* BEL="X29/Y12/lc6" *)
   SB_DFF  dff_29_94 (
      .C       (i_clk         ),
      .D       (p2_dl[94]    ),
      .Q       (p3_dl[94]    )
   );
   (* BEL="X2/Y12/lc7" *)
   SB_DFF  dff_2_95 (
      .C       (i_clk         ),
      .D       (p0_dl[96]  ),
      .Q       (p1_dl[95]    )
   );

   (* BEL="X3/Y12/lc7" *)
   SB_DFF  dff_3_95 (
      .C       (i_clk         ),
      .D       (p1_dl[95]    ),
      .Q       (p2_dl[95]    )
   );


   (* BEL="X29/Y12/lc7" *)
   SB_DFF  dff_29_95 (
      .C       (i_clk         ),
      .D       (p2_dl[95]    ),
      .Q       (p3_dl[95]    )
   );
   (* BEL="X2/Y13/lc0" *)
   SB_DFF  dff_2_96 (
      .C       (i_clk         ),
      .D       (p0_dl[97]  ),
      .Q       (p1_dl[96]    )
   );

   (* BEL="X3/Y13/lc0" *)
   SB_DFF  dff_3_96 (
      .C       (i_clk         ),
      .D       (p1_dl[96]    ),
      .Q       (p2_dl[96]    )
   );


   (* BEL="X29/Y13/lc0" *)
   SB_DFF  dff_29_96 (
      .C       (i_clk         ),
      .D       (p2_dl[96]    ),
      .Q       (p3_dl[96]    )
   );
   (* BEL="X2/Y13/lc1" *)
   SB_DFF  dff_2_97 (
      .C       (i_clk         ),
      .D       (p0_dl[98]  ),
      .Q       (p1_dl[97]    )
   );

   (* BEL="X3/Y13/lc1" *)
   SB_DFF  dff_3_97 (
      .C       (i_clk         ),
      .D       (p1_dl[97]    ),
      .Q       (p2_dl[97]    )
   );


   (* BEL="X29/Y13/lc1" *)
   SB_DFF  dff_29_97 (
      .C       (i_clk         ),
      .D       (p2_dl[97]    ),
      .Q       (p3_dl[97]    )
   );
   (* BEL="X2/Y13/lc2" *)
   SB_DFF  dff_2_98 (
      .C       (i_clk         ),
      .D       (p0_dl[99]  ),
      .Q       (p1_dl[98]    )
   );

   (* BEL="X3/Y13/lc2" *)
   SB_DFF  dff_3_98 (
      .C       (i_clk         ),
      .D       (p1_dl[98]    ),
      .Q       (p2_dl[98]    )
   );


   (* BEL="X29/Y13/lc2" *)
   SB_DFF  dff_29_98 (
      .C       (i_clk         ),
      .D       (p2_dl[98]    ),
      .Q       (p3_dl[98]    )
   );
   (* BEL="X2/Y13/lc3" *)
   SB_DFF  dff_2_99 (
      .C       (i_clk         ),
      .D       (p0_dl[100]  ),
      .Q       (p1_dl[99]    )
   );

   (* BEL="X3/Y13/lc3" *)
   SB_DFF  dff_3_99 (
      .C       (i_clk         ),
      .D       (p1_dl[99]    ),
      .Q       (p2_dl[99]    )
   );


   (* BEL="X29/Y13/lc3" *)
   SB_DFF  dff_29_99 (
      .C       (i_clk         ),
      .D       (p2_dl[99]    ),
      .Q       (p3_dl[99]    )
   );
   (* BEL="X2/Y13/lc4" *)
   SB_DFF  dff_2_100 (
      .C       (i_clk         ),
      .D       (p0_dl[101]  ),
      .Q       (p1_dl[100]    )
   );

   (* BEL="X3/Y13/lc4" *)
   SB_DFF  dff_3_100 (
      .C       (i_clk         ),
      .D       (p1_dl[100]    ),
      .Q       (p2_dl[100]    )
   );


   (* BEL="X29/Y13/lc4" *)
   SB_DFF  dff_29_100 (
      .C       (i_clk         ),
      .D       (p2_dl[100]    ),
      .Q       (p3_dl[100]    )
   );
   (* BEL="X2/Y13/lc5" *)
   SB_DFF  dff_2_101 (
      .C       (i_clk         ),
      .D       (p0_dl[102]  ),
      .Q       (p1_dl[101]    )
   );

   (* BEL="X3/Y13/lc5" *)
   SB_DFF  dff_3_101 (
      .C       (i_clk         ),
      .D       (p1_dl[101]    ),
      .Q       (p2_dl[101]    )
   );


   (* BEL="X29/Y13/lc5" *)
   SB_DFF  dff_29_101 (
      .C       (i_clk         ),
      .D       (p2_dl[101]    ),
      .Q       (p3_dl[101]    )
   );
   (* BEL="X2/Y13/lc6" *)
   SB_DFF  dff_2_102 (
      .C       (i_clk         ),
      .D       (p0_dl[103]  ),
      .Q       (p1_dl[102]    )
   );

   (* BEL="X3/Y13/lc6" *)
   SB_DFF  dff_3_102 (
      .C       (i_clk         ),
      .D       (p1_dl[102]    ),
      .Q       (p2_dl[102]    )
   );


   (* BEL="X29/Y13/lc6" *)
   SB_DFF  dff_29_102 (
      .C       (i_clk         ),
      .D       (p2_dl[102]    ),
      .Q       (p3_dl[102]    )
   );
   (* BEL="X2/Y13/lc7" *)
   SB_DFF  dff_2_103 (
      .C       (i_clk         ),
      .D       (p0_dl[104]  ),
      .Q       (p1_dl[103]    )
   );

   (* BEL="X3/Y13/lc7" *)
   SB_DFF  dff_3_103 (
      .C       (i_clk         ),
      .D       (p1_dl[103]    ),
      .Q       (p2_dl[103]    )
   );


   (* BEL="X29/Y13/lc7" *)
   SB_DFF  dff_29_103 (
      .C       (i_clk         ),
      .D       (p2_dl[103]    ),
      .Q       (p3_dl[103]    )
   );
   (* BEL="X2/Y14/lc0" *)
   SB_DFF  dff_2_104 (
      .C       (i_clk         ),
      .D       (p0_dl[105]  ),
      .Q       (p1_dl[104]    )
   );

   (* BEL="X3/Y14/lc0" *)
   SB_DFF  dff_3_104 (
      .C       (i_clk         ),
      .D       (p1_dl[104]    ),
      .Q       (p2_dl[104]    )
   );


   (* BEL="X29/Y14/lc0" *)
   SB_DFF  dff_29_104 (
      .C       (i_clk         ),
      .D       (p2_dl[104]    ),
      .Q       (p3_dl[104]    )
   );
   (* BEL="X2/Y14/lc1" *)
   SB_DFF  dff_2_105 (
      .C       (i_clk         ),
      .D       (p0_dl[106]  ),
      .Q       (p1_dl[105]    )
   );

   (* BEL="X3/Y14/lc1" *)
   SB_DFF  dff_3_105 (
      .C       (i_clk         ),
      .D       (p1_dl[105]    ),
      .Q       (p2_dl[105]    )
   );


   (* BEL="X29/Y14/lc1" *)
   SB_DFF  dff_29_105 (
      .C       (i_clk         ),
      .D       (p2_dl[105]    ),
      .Q       (p3_dl[105]    )
   );
   (* BEL="X2/Y14/lc2" *)
   SB_DFF  dff_2_106 (
      .C       (i_clk         ),
      .D       (p0_dl[107]  ),
      .Q       (p1_dl[106]    )
   );

   (* BEL="X3/Y14/lc2" *)
   SB_DFF  dff_3_106 (
      .C       (i_clk         ),
      .D       (p1_dl[106]    ),
      .Q       (p2_dl[106]    )
   );


   (* BEL="X29/Y14/lc2" *)
   SB_DFF  dff_29_106 (
      .C       (i_clk         ),
      .D       (p2_dl[106]    ),
      .Q       (p3_dl[106]    )
   );
   (* BEL="X2/Y14/lc3" *)
   SB_DFF  dff_2_107 (
      .C       (i_clk         ),
      .D       (p0_dl[108]  ),
      .Q       (p1_dl[107]    )
   );

   (* BEL="X3/Y14/lc3" *)
   SB_DFF  dff_3_107 (
      .C       (i_clk         ),
      .D       (p1_dl[107]    ),
      .Q       (p2_dl[107]    )
   );


   (* BEL="X29/Y14/lc3" *)
   SB_DFF  dff_29_107 (
      .C       (i_clk         ),
      .D       (p2_dl[107]    ),
      .Q       (p3_dl[107]    )
   );
   (* BEL="X2/Y14/lc4" *)
   SB_DFF  dff_2_108 (
      .C       (i_clk         ),
      .D       (p0_dl[109]  ),
      .Q       (p1_dl[108]    )
   );

   (* BEL="X3/Y14/lc4" *)
   SB_DFF  dff_3_108 (
      .C       (i_clk         ),
      .D       (p1_dl[108]    ),
      .Q       (p2_dl[108]    )
   );


   (* BEL="X29/Y14/lc4" *)
   SB_DFF  dff_29_108 (
      .C       (i_clk         ),
      .D       (p2_dl[108]    ),
      .Q       (p3_dl[108]    )
   );
   (* BEL="X2/Y14/lc5" *)
   SB_DFF  dff_2_109 (
      .C       (i_clk         ),
      .D       (p0_dl[110]  ),
      .Q       (p1_dl[109]    )
   );

   (* BEL="X3/Y14/lc5" *)
   SB_DFF  dff_3_109 (
      .C       (i_clk         ),
      .D       (p1_dl[109]    ),
      .Q       (p2_dl[109]    )
   );


   (* BEL="X29/Y14/lc5" *)
   SB_DFF  dff_29_109 (
      .C       (i_clk         ),
      .D       (p2_dl[109]    ),
      .Q       (p3_dl[109]    )
   );
   (* BEL="X2/Y14/lc6" *)
   SB_DFF  dff_2_110 (
      .C       (i_clk         ),
      .D       (p0_dl[111]  ),
      .Q       (p1_dl[110]    )
   );

   (* BEL="X3/Y14/lc6" *)
   SB_DFF  dff_3_110 (
      .C       (i_clk         ),
      .D       (p1_dl[110]    ),
      .Q       (p2_dl[110]    )
   );


   (* BEL="X29/Y14/lc6" *)
   SB_DFF  dff_29_110 (
      .C       (i_clk         ),
      .D       (p2_dl[110]    ),
      .Q       (p3_dl[110]    )
   );
   (* BEL="X2/Y14/lc7" *)
   SB_DFF  dff_2_111 (
      .C       (i_clk         ),
      .D       (p0_dl[112]  ),
      .Q       (p1_dl[111]    )
   );

   (* BEL="X3/Y14/lc7" *)
   SB_DFF  dff_3_111 (
      .C       (i_clk         ),
      .D       (p1_dl[111]    ),
      .Q       (p2_dl[111]    )
   );


   (* BEL="X29/Y14/lc7" *)
   SB_DFF  dff_29_111 (
      .C       (i_clk         ),
      .D       (p2_dl[111]    ),
      .Q       (p3_dl[111]    )
   );
   (* BEL="X2/Y15/lc0" *)
   SB_DFF  dff_2_112 (
      .C       (i_clk         ),
      .D       (p0_dl[113]  ),
      .Q       (p1_dl[112]    )
   );

   (* BEL="X3/Y15/lc0" *)
   SB_DFF  dff_3_112 (
      .C       (i_clk         ),
      .D       (p1_dl[112]    ),
      .Q       (p2_dl[112]    )
   );


   (* BEL="X29/Y15/lc0" *)
   SB_DFF  dff_29_112 (
      .C       (i_clk         ),
      .D       (p2_dl[112]    ),
      .Q       (p3_dl[112]    )
   );
   (* BEL="X2/Y15/lc1" *)
   SB_DFF  dff_2_113 (
      .C       (i_clk         ),
      .D       (p0_dl[114]  ),
      .Q       (p1_dl[113]    )
   );

   (* BEL="X3/Y15/lc1" *)
   SB_DFF  dff_3_113 (
      .C       (i_clk         ),
      .D       (p1_dl[113]    ),
      .Q       (p2_dl[113]    )
   );


   (* BEL="X29/Y15/lc1" *)
   SB_DFF  dff_29_113 (
      .C       (i_clk         ),
      .D       (p2_dl[113]    ),
      .Q       (p3_dl[113]    )
   );
   (* BEL="X2/Y15/lc2" *)
   SB_DFF  dff_2_114 (
      .C       (i_clk         ),
      .D       (p0_dl[115]  ),
      .Q       (p1_dl[114]    )
   );

   (* BEL="X3/Y15/lc2" *)
   SB_DFF  dff_3_114 (
      .C       (i_clk         ),
      .D       (p1_dl[114]    ),
      .Q       (p2_dl[114]    )
   );


   (* BEL="X29/Y15/lc2" *)
   SB_DFF  dff_29_114 (
      .C       (i_clk         ),
      .D       (p2_dl[114]    ),
      .Q       (p3_dl[114]    )
   );
   (* BEL="X2/Y15/lc3" *)
   SB_DFF  dff_2_115 (
      .C       (i_clk         ),
      .D       (p0_dl[116]  ),
      .Q       (p1_dl[115]    )
   );

   (* BEL="X3/Y15/lc3" *)
   SB_DFF  dff_3_115 (
      .C       (i_clk         ),
      .D       (p1_dl[115]    ),
      .Q       (p2_dl[115]    )
   );


   (* BEL="X29/Y15/lc3" *)
   SB_DFF  dff_29_115 (
      .C       (i_clk         ),
      .D       (p2_dl[115]    ),
      .Q       (p3_dl[115]    )
   );
   (* BEL="X2/Y15/lc4" *)
   SB_DFF  dff_2_116 (
      .C       (i_clk         ),
      .D       (p0_dl[117]  ),
      .Q       (p1_dl[116]    )
   );

   (* BEL="X3/Y15/lc4" *)
   SB_DFF  dff_3_116 (
      .C       (i_clk         ),
      .D       (p1_dl[116]    ),
      .Q       (p2_dl[116]    )
   );


   (* BEL="X29/Y15/lc4" *)
   SB_DFF  dff_29_116 (
      .C       (i_clk         ),
      .D       (p2_dl[116]    ),
      .Q       (p3_dl[116]    )
   );
   (* BEL="X2/Y15/lc5" *)
   SB_DFF  dff_2_117 (
      .C       (i_clk         ),
      .D       (p0_dl[118]  ),
      .Q       (p1_dl[117]    )
   );

   (* BEL="X3/Y15/lc5" *)
   SB_DFF  dff_3_117 (
      .C       (i_clk         ),
      .D       (p1_dl[117]    ),
      .Q       (p2_dl[117]    )
   );


   (* BEL="X29/Y15/lc5" *)
   SB_DFF  dff_29_117 (
      .C       (i_clk         ),
      .D       (p2_dl[117]    ),
      .Q       (p3_dl[117]    )
   );
   (* BEL="X2/Y15/lc6" *)
   SB_DFF  dff_2_118 (
      .C       (i_clk         ),
      .D       (p0_dl[119]  ),
      .Q       (p1_dl[118]    )
   );

   (* BEL="X3/Y15/lc6" *)
   SB_DFF  dff_3_118 (
      .C       (i_clk         ),
      .D       (p1_dl[118]    ),
      .Q       (p2_dl[118]    )
   );


   (* BEL="X29/Y15/lc6" *)
   SB_DFF  dff_29_118 (
      .C       (i_clk         ),
      .D       (p2_dl[118]    ),
      .Q       (p3_dl[118]    )
   );
   (* BEL="X2/Y15/lc7" *)
   SB_DFF  dff_2_119 (
      .C       (i_clk         ),
      .D       (p0_dl[120]  ),
      .Q       (p1_dl[119]    )
   );

   (* BEL="X3/Y15/lc7" *)
   SB_DFF  dff_3_119 (
      .C       (i_clk         ),
      .D       (p1_dl[119]    ),
      .Q       (p2_dl[119]    )
   );


   (* BEL="X29/Y15/lc7" *)
   SB_DFF  dff_29_119 (
      .C       (i_clk         ),
      .D       (p2_dl[119]    ),
      .Q       (p3_dl[119]    )
   );
   (* BEL="X2/Y16/lc0" *)
   SB_DFF  dff_2_120 (
      .C       (i_clk         ),
      .D       (p0_dl[121]  ),
      .Q       (p1_dl[120]    )
   );

   (* BEL="X3/Y16/lc0" *)
   SB_DFF  dff_3_120 (
      .C       (i_clk         ),
      .D       (p1_dl[120]    ),
      .Q       (p2_dl[120]    )
   );


   (* BEL="X29/Y16/lc0" *)
   SB_DFF  dff_29_120 (
      .C       (i_clk         ),
      .D       (p2_dl[120]    ),
      .Q       (p3_dl[120]    )
   );
   (* BEL="X2/Y16/lc1" *)
   SB_DFF  dff_2_121 (
      .C       (i_clk         ),
      .D       (p0_dl[122]  ),
      .Q       (p1_dl[121]    )
   );

   (* BEL="X3/Y16/lc1" *)
   SB_DFF  dff_3_121 (
      .C       (i_clk         ),
      .D       (p1_dl[121]    ),
      .Q       (p2_dl[121]    )
   );


   (* BEL="X29/Y16/lc1" *)
   SB_DFF  dff_29_121 (
      .C       (i_clk         ),
      .D       (p2_dl[121]    ),
      .Q       (p3_dl[121]    )
   );
   (* BEL="X2/Y16/lc2" *)
   SB_DFF  dff_2_122 (
      .C       (i_clk         ),
      .D       (p0_dl[123]  ),
      .Q       (p1_dl[122]    )
   );

   (* BEL="X3/Y16/lc2" *)
   SB_DFF  dff_3_122 (
      .C       (i_clk         ),
      .D       (p1_dl[122]    ),
      .Q       (p2_dl[122]    )
   );


   (* BEL="X29/Y16/lc2" *)
   SB_DFF  dff_29_122 (
      .C       (i_clk         ),
      .D       (p2_dl[122]    ),
      .Q       (p3_dl[122]    )
   );
   (* BEL="X2/Y16/lc3" *)
   SB_DFF  dff_2_123 (
      .C       (i_clk         ),
      .D       (p0_dl[124]  ),
      .Q       (p1_dl[123]    )
   );

   (* BEL="X3/Y16/lc3" *)
   SB_DFF  dff_3_123 (
      .C       (i_clk         ),
      .D       (p1_dl[123]    ),
      .Q       (p2_dl[123]    )
   );


   (* BEL="X29/Y16/lc3" *)
   SB_DFF  dff_29_123 (
      .C       (i_clk         ),
      .D       (p2_dl[123]    ),
      .Q       (p3_dl[123]    )
   );
   (* BEL="X2/Y16/lc4" *)
   SB_DFF  dff_2_124 (
      .C       (i_clk         ),
      .D       (p0_dl[125]  ),
      .Q       (p1_dl[124]    )
   );

   (* BEL="X3/Y16/lc4" *)
   SB_DFF  dff_3_124 (
      .C       (i_clk         ),
      .D       (p1_dl[124]    ),
      .Q       (p2_dl[124]    )
   );


   (* BEL="X29/Y16/lc4" *)
   SB_DFF  dff_29_124 (
      .C       (i_clk         ),
      .D       (p2_dl[124]    ),
      .Q       (p3_dl[124]    )
   );
   (* BEL="X2/Y16/lc5" *)
   SB_DFF  dff_2_125 (
      .C       (i_clk         ),
      .D       (p0_dl[126]  ),
      .Q       (p1_dl[125]    )
   );

   (* BEL="X3/Y16/lc5" *)
   SB_DFF  dff_3_125 (
      .C       (i_clk         ),
      .D       (p1_dl[125]    ),
      .Q       (p2_dl[125]    )
   );


   (* BEL="X29/Y16/lc5" *)
   SB_DFF  dff_29_125 (
      .C       (i_clk         ),
      .D       (p2_dl[125]    ),
      .Q       (p3_dl[125]    )
   );
   (* BEL="X2/Y16/lc6" *)
   SB_DFF  dff_2_126 (
      .C       (i_clk         ),
      .D       (p0_dl[127]  ),
      .Q       (p1_dl[126]    )
   );

   (* BEL="X3/Y16/lc6" *)
   SB_DFF  dff_3_126 (
      .C       (i_clk         ),
      .D       (p1_dl[126]    ),
      .Q       (p2_dl[126]    )
   );


   (* BEL="X29/Y16/lc6" *)
   SB_DFF  dff_29_126 (
      .C       (i_clk         ),
      .D       (p2_dl[126]    ),
      .Q       (p3_dl[126]    )
   );
   (* BEL="X2/Y16/lc7" *)
   SB_DFF  dff_2_127 (
      .C       (i_clk         ),
      .D       (p0_dl[128]  ),
      .Q       (p1_dl[127]    )
   );

   (* BEL="X3/Y16/lc7" *)
   SB_DFF  dff_3_127 (
      .C       (i_clk         ),
      .D       (p1_dl[127]    ),
      .Q       (p2_dl[127]    )
   );


   (* BEL="X29/Y16/lc7" *)
   SB_DFF  dff_29_127 (
      .C       (i_clk         ),
      .D       (p2_dl[127]    ),
      .Q       (p3_dl[127]    )
   );
   (* BEL="X2/Y17/lc0" *)
   SB_DFF  dff_2_128 (
      .C       (i_clk         ),
      .D       (p0_dl[129]  ),
      .Q       (p1_dl[128]    )
   );

   (* BEL="X3/Y17/lc0" *)
   SB_DFF  dff_3_128 (
      .C       (i_clk         ),
      .D       (p1_dl[128]    ),
      .Q       (p2_dl[128]    )
   );


   (* BEL="X29/Y17/lc0" *)
   SB_DFF  dff_29_128 (
      .C       (i_clk         ),
      .D       (p2_dl[128]    ),
      .Q       (p3_dl[128]    )
   );
   (* BEL="X2/Y17/lc1" *)
   SB_DFF  dff_2_129 (
      .C       (i_clk         ),
      .D       (p0_dl[130]  ),
      .Q       (p1_dl[129]    )
   );

   (* BEL="X3/Y17/lc1" *)
   SB_DFF  dff_3_129 (
      .C       (i_clk         ),
      .D       (p1_dl[129]    ),
      .Q       (p2_dl[129]    )
   );


   (* BEL="X29/Y17/lc1" *)
   SB_DFF  dff_29_129 (
      .C       (i_clk         ),
      .D       (p2_dl[129]    ),
      .Q       (p3_dl[129]    )
   );
   (* BEL="X2/Y17/lc2" *)
   SB_DFF  dff_2_130 (
      .C       (i_clk         ),
      .D       (p0_dl[131]  ),
      .Q       (p1_dl[130]    )
   );

   (* BEL="X3/Y17/lc2" *)
   SB_DFF  dff_3_130 (
      .C       (i_clk         ),
      .D       (p1_dl[130]    ),
      .Q       (p2_dl[130]    )
   );


   (* BEL="X29/Y17/lc2" *)
   SB_DFF  dff_29_130 (
      .C       (i_clk         ),
      .D       (p2_dl[130]    ),
      .Q       (p3_dl[130]    )
   );
   (* BEL="X2/Y17/lc3" *)
   SB_DFF  dff_2_131 (
      .C       (i_clk         ),
      .D       (p0_dl[132]  ),
      .Q       (p1_dl[131]    )
   );

   (* BEL="X3/Y17/lc3" *)
   SB_DFF  dff_3_131 (
      .C       (i_clk         ),
      .D       (p1_dl[131]    ),
      .Q       (p2_dl[131]    )
   );


   (* BEL="X29/Y17/lc3" *)
   SB_DFF  dff_29_131 (
      .C       (i_clk         ),
      .D       (p2_dl[131]    ),
      .Q       (p3_dl[131]    )
   );
   (* BEL="X2/Y17/lc4" *)
   SB_DFF  dff_2_132 (
      .C       (i_clk         ),
      .D       (p0_dl[133]  ),
      .Q       (p1_dl[132]    )
   );

   (* BEL="X3/Y17/lc4" *)
   SB_DFF  dff_3_132 (
      .C       (i_clk         ),
      .D       (p1_dl[132]    ),
      .Q       (p2_dl[132]    )
   );


   (* BEL="X29/Y17/lc4" *)
   SB_DFF  dff_29_132 (
      .C       (i_clk         ),
      .D       (p2_dl[132]    ),
      .Q       (p3_dl[132]    )
   );
   (* BEL="X2/Y17/lc5" *)
   SB_DFF  dff_2_133 (
      .C       (i_clk         ),
      .D       (p0_dl[134]  ),
      .Q       (p1_dl[133]    )
   );

   (* BEL="X3/Y17/lc5" *)
   SB_DFF  dff_3_133 (
      .C       (i_clk         ),
      .D       (p1_dl[133]    ),
      .Q       (p2_dl[133]    )
   );


   (* BEL="X29/Y17/lc5" *)
   SB_DFF  dff_29_133 (
      .C       (i_clk         ),
      .D       (p2_dl[133]    ),
      .Q       (p3_dl[133]    )
   );
   (* BEL="X2/Y17/lc6" *)
   SB_DFF  dff_2_134 (
      .C       (i_clk         ),
      .D       (p0_dl[135]  ),
      .Q       (p1_dl[134]    )
   );

   (* BEL="X3/Y17/lc6" *)
   SB_DFF  dff_3_134 (
      .C       (i_clk         ),
      .D       (p1_dl[134]    ),
      .Q       (p2_dl[134]    )
   );


   (* BEL="X29/Y17/lc6" *)
   SB_DFF  dff_29_134 (
      .C       (i_clk         ),
      .D       (p2_dl[134]    ),
      .Q       (p3_dl[134]    )
   );
   (* BEL="X2/Y17/lc7" *)
   SB_DFF  dff_2_135 (
      .C       (i_clk         ),
      .D       (p0_dl[136]  ),
      .Q       (p1_dl[135]    )
   );

   (* BEL="X3/Y17/lc7" *)
   SB_DFF  dff_3_135 (
      .C       (i_clk         ),
      .D       (p1_dl[135]    ),
      .Q       (p2_dl[135]    )
   );


   (* BEL="X29/Y17/lc7" *)
   SB_DFF  dff_29_135 (
      .C       (i_clk         ),
      .D       (p2_dl[135]    ),
      .Q       (p3_dl[135]    )
   );
   (* BEL="X2/Y18/lc0" *)
   SB_DFF  dff_2_136 (
      .C       (i_clk         ),
      .D       (p0_dl[137]  ),
      .Q       (p1_dl[136]    )
   );

   (* BEL="X3/Y18/lc0" *)
   SB_DFF  dff_3_136 (
      .C       (i_clk         ),
      .D       (p1_dl[136]    ),
      .Q       (p2_dl[136]    )
   );


   (* BEL="X29/Y18/lc0" *)
   SB_DFF  dff_29_136 (
      .C       (i_clk         ),
      .D       (p2_dl[136]    ),
      .Q       (p3_dl[136]    )
   );
   (* BEL="X2/Y18/lc1" *)
   SB_DFF  dff_2_137 (
      .C       (i_clk         ),
      .D       (p0_dl[138]  ),
      .Q       (p1_dl[137]    )
   );

   (* BEL="X3/Y18/lc1" *)
   SB_DFF  dff_3_137 (
      .C       (i_clk         ),
      .D       (p1_dl[137]    ),
      .Q       (p2_dl[137]    )
   );


   (* BEL="X29/Y18/lc1" *)
   SB_DFF  dff_29_137 (
      .C       (i_clk         ),
      .D       (p2_dl[137]    ),
      .Q       (p3_dl[137]    )
   );
   (* BEL="X2/Y18/lc2" *)
   SB_DFF  dff_2_138 (
      .C       (i_clk         ),
      .D       (p0_dl[139]  ),
      .Q       (p1_dl[138]    )
   );

   (* BEL="X3/Y18/lc2" *)
   SB_DFF  dff_3_138 (
      .C       (i_clk         ),
      .D       (p1_dl[138]    ),
      .Q       (p2_dl[138]    )
   );


   (* BEL="X29/Y18/lc2" *)
   SB_DFF  dff_29_138 (
      .C       (i_clk         ),
      .D       (p2_dl[138]    ),
      .Q       (p3_dl[138]    )
   );
   (* BEL="X2/Y18/lc3" *)
   SB_DFF  dff_2_139 (
      .C       (i_clk         ),
      .D       (p0_dl[140]  ),
      .Q       (p1_dl[139]    )
   );

   (* BEL="X3/Y18/lc3" *)
   SB_DFF  dff_3_139 (
      .C       (i_clk         ),
      .D       (p1_dl[139]    ),
      .Q       (p2_dl[139]    )
   );


   (* BEL="X29/Y18/lc3" *)
   SB_DFF  dff_29_139 (
      .C       (i_clk         ),
      .D       (p2_dl[139]    ),
      .Q       (p3_dl[139]    )
   );
   (* BEL="X2/Y18/lc4" *)
   SB_DFF  dff_2_140 (
      .C       (i_clk         ),
      .D       (p0_dl[141]  ),
      .Q       (p1_dl[140]    )
   );

   (* BEL="X3/Y18/lc4" *)
   SB_DFF  dff_3_140 (
      .C       (i_clk         ),
      .D       (p1_dl[140]    ),
      .Q       (p2_dl[140]    )
   );


   (* BEL="X29/Y18/lc4" *)
   SB_DFF  dff_29_140 (
      .C       (i_clk         ),
      .D       (p2_dl[140]    ),
      .Q       (p3_dl[140]    )
   );
   (* BEL="X2/Y18/lc5" *)
   SB_DFF  dff_2_141 (
      .C       (i_clk         ),
      .D       (p0_dl[142]  ),
      .Q       (p1_dl[141]    )
   );

   (* BEL="X3/Y18/lc5" *)
   SB_DFF  dff_3_141 (
      .C       (i_clk         ),
      .D       (p1_dl[141]    ),
      .Q       (p2_dl[141]    )
   );


   (* BEL="X29/Y18/lc5" *)
   SB_DFF  dff_29_141 (
      .C       (i_clk         ),
      .D       (p2_dl[141]    ),
      .Q       (p3_dl[141]    )
   );
   (* BEL="X2/Y18/lc6" *)
   SB_DFF  dff_2_142 (
      .C       (i_clk         ),
      .D       (p0_dl[143]  ),
      .Q       (p1_dl[142]    )
   );

   (* BEL="X3/Y18/lc6" *)
   SB_DFF  dff_3_142 (
      .C       (i_clk         ),
      .D       (p1_dl[142]    ),
      .Q       (p2_dl[142]    )
   );


   (* BEL="X29/Y18/lc6" *)
   SB_DFF  dff_29_142 (
      .C       (i_clk         ),
      .D       (p2_dl[142]    ),
      .Q       (p3_dl[142]    )
   );
   (* BEL="X2/Y18/lc7" *)
   SB_DFF  dff_2_143 (
      .C       (i_clk         ),
      .D       (p0_dl[144]  ),
      .Q       (p1_dl[143]    )
   );

   (* BEL="X3/Y18/lc7" *)
   SB_DFF  dff_3_143 (
      .C       (i_clk         ),
      .D       (p1_dl[143]    ),
      .Q       (p2_dl[143]    )
   );


   (* BEL="X29/Y18/lc7" *)
   SB_DFF  dff_29_143 (
      .C       (i_clk         ),
      .D       (p2_dl[143]    ),
      .Q       (p3_dl[143]    )
   );
   (* BEL="X2/Y19/lc0" *)
   SB_DFF  dff_2_144 (
      .C       (i_clk         ),
      .D       (p0_dl[145]  ),
      .Q       (p1_dl[144]    )
   );

   (* BEL="X3/Y19/lc0" *)
   SB_DFF  dff_3_144 (
      .C       (i_clk         ),
      .D       (p1_dl[144]    ),
      .Q       (p2_dl[144]    )
   );


   (* BEL="X29/Y19/lc0" *)
   SB_DFF  dff_29_144 (
      .C       (i_clk         ),
      .D       (p2_dl[144]    ),
      .Q       (p3_dl[144]    )
   );
   (* BEL="X2/Y19/lc1" *)
   SB_DFF  dff_2_145 (
      .C       (i_clk         ),
      .D       (p0_dl[146]  ),
      .Q       (p1_dl[145]    )
   );

   (* BEL="X3/Y19/lc1" *)
   SB_DFF  dff_3_145 (
      .C       (i_clk         ),
      .D       (p1_dl[145]    ),
      .Q       (p2_dl[145]    )
   );


   (* BEL="X29/Y19/lc1" *)
   SB_DFF  dff_29_145 (
      .C       (i_clk         ),
      .D       (p2_dl[145]    ),
      .Q       (p3_dl[145]    )
   );
   (* BEL="X2/Y19/lc2" *)
   SB_DFF  dff_2_146 (
      .C       (i_clk         ),
      .D       (p0_dl[147]  ),
      .Q       (p1_dl[146]    )
   );

   (* BEL="X3/Y19/lc2" *)
   SB_DFF  dff_3_146 (
      .C       (i_clk         ),
      .D       (p1_dl[146]    ),
      .Q       (p2_dl[146]    )
   );


   (* BEL="X29/Y19/lc2" *)
   SB_DFF  dff_29_146 (
      .C       (i_clk         ),
      .D       (p2_dl[146]    ),
      .Q       (p3_dl[146]    )
   );
   (* BEL="X2/Y19/lc3" *)
   SB_DFF  dff_2_147 (
      .C       (i_clk         ),
      .D       (p0_dl[148]  ),
      .Q       (p1_dl[147]    )
   );

   (* BEL="X3/Y19/lc3" *)
   SB_DFF  dff_3_147 (
      .C       (i_clk         ),
      .D       (p1_dl[147]    ),
      .Q       (p2_dl[147]    )
   );


   (* BEL="X29/Y19/lc3" *)
   SB_DFF  dff_29_147 (
      .C       (i_clk         ),
      .D       (p2_dl[147]    ),
      .Q       (p3_dl[147]    )
   );
   (* BEL="X2/Y19/lc4" *)
   SB_DFF  dff_2_148 (
      .C       (i_clk         ),
      .D       (p0_dl[149]  ),
      .Q       (p1_dl[148]    )
   );

   (* BEL="X3/Y19/lc4" *)
   SB_DFF  dff_3_148 (
      .C       (i_clk         ),
      .D       (p1_dl[148]    ),
      .Q       (p2_dl[148]    )
   );


   (* BEL="X29/Y19/lc4" *)
   SB_DFF  dff_29_148 (
      .C       (i_clk         ),
      .D       (p2_dl[148]    ),
      .Q       (p3_dl[148]    )
   );
   (* BEL="X2/Y19/lc5" *)
   SB_DFF  dff_2_149 (
      .C       (i_clk         ),
      .D       (p0_dl[150]  ),
      .Q       (p1_dl[149]    )
   );

   (* BEL="X3/Y19/lc5" *)
   SB_DFF  dff_3_149 (
      .C       (i_clk         ),
      .D       (p1_dl[149]    ),
      .Q       (p2_dl[149]    )
   );


   (* BEL="X29/Y19/lc5" *)
   SB_DFF  dff_29_149 (
      .C       (i_clk         ),
      .D       (p2_dl[149]    ),
      .Q       (p3_dl[149]    )
   );
   (* BEL="X2/Y19/lc6" *)
   SB_DFF  dff_2_150 (
      .C       (i_clk         ),
      .D       (p0_dl[151]  ),
      .Q       (p1_dl[150]    )
   );

   (* BEL="X3/Y19/lc6" *)
   SB_DFF  dff_3_150 (
      .C       (i_clk         ),
      .D       (p1_dl[150]    ),
      .Q       (p2_dl[150]    )
   );


   (* BEL="X29/Y19/lc6" *)
   SB_DFF  dff_29_150 (
      .C       (i_clk         ),
      .D       (p2_dl[150]    ),
      .Q       (p3_dl[150]    )
   );
   (* BEL="X2/Y19/lc7" *)
   SB_DFF  dff_2_151 (
      .C       (i_clk         ),
      .D       (p0_dl[152]  ),
      .Q       (p1_dl[151]    )
   );

   (* BEL="X3/Y19/lc7" *)
   SB_DFF  dff_3_151 (
      .C       (i_clk         ),
      .D       (p1_dl[151]    ),
      .Q       (p2_dl[151]    )
   );


   (* BEL="X29/Y19/lc7" *)
   SB_DFF  dff_29_151 (
      .C       (i_clk         ),
      .D       (p2_dl[151]    ),
      .Q       (p3_dl[151]    )
   );
   (* BEL="X2/Y20/lc0" *)
   SB_DFF  dff_2_152 (
      .C       (i_clk         ),
      .D       (p0_dl[153]  ),
      .Q       (p1_dl[152]    )
   );

   (* BEL="X3/Y20/lc0" *)
   SB_DFF  dff_3_152 (
      .C       (i_clk         ),
      .D       (p1_dl[152]    ),
      .Q       (p2_dl[152]    )
   );


   (* BEL="X29/Y20/lc0" *)
   SB_DFF  dff_29_152 (
      .C       (i_clk         ),
      .D       (p2_dl[152]    ),
      .Q       (p3_dl[152]    )
   );
   (* BEL="X2/Y20/lc1" *)
   SB_DFF  dff_2_153 (
      .C       (i_clk         ),
      .D       (p0_dl[154]  ),
      .Q       (p1_dl[153]    )
   );

   (* BEL="X3/Y20/lc1" *)
   SB_DFF  dff_3_153 (
      .C       (i_clk         ),
      .D       (p1_dl[153]    ),
      .Q       (p2_dl[153]    )
   );


   (* BEL="X29/Y20/lc1" *)
   SB_DFF  dff_29_153 (
      .C       (i_clk         ),
      .D       (p2_dl[153]    ),
      .Q       (p3_dl[153]    )
   );
   (* BEL="X2/Y20/lc2" *)
   SB_DFF  dff_2_154 (
      .C       (i_clk         ),
      .D       (p0_dl[155]  ),
      .Q       (p1_dl[154]    )
   );

   (* BEL="X3/Y20/lc2" *)
   SB_DFF  dff_3_154 (
      .C       (i_clk         ),
      .D       (p1_dl[154]    ),
      .Q       (p2_dl[154]    )
   );


   (* BEL="X29/Y20/lc2" *)
   SB_DFF  dff_29_154 (
      .C       (i_clk         ),
      .D       (p2_dl[154]    ),
      .Q       (p3_dl[154]    )
   );
   (* BEL="X2/Y20/lc3" *)
   SB_DFF  dff_2_155 (
      .C       (i_clk         ),
      .D       (p0_dl[156]  ),
      .Q       (p1_dl[155]    )
   );

   (* BEL="X3/Y20/lc3" *)
   SB_DFF  dff_3_155 (
      .C       (i_clk         ),
      .D       (p1_dl[155]    ),
      .Q       (p2_dl[155]    )
   );


   (* BEL="X29/Y20/lc3" *)
   SB_DFF  dff_29_155 (
      .C       (i_clk         ),
      .D       (p2_dl[155]    ),
      .Q       (p3_dl[155]    )
   );
   (* BEL="X2/Y20/lc4" *)
   SB_DFF  dff_2_156 (
      .C       (i_clk         ),
      .D       (p0_dl[157]  ),
      .Q       (p1_dl[156]    )
   );

   (* BEL="X3/Y20/lc4" *)
   SB_DFF  dff_3_156 (
      .C       (i_clk         ),
      .D       (p1_dl[156]    ),
      .Q       (p2_dl[156]    )
   );


   (* BEL="X29/Y20/lc4" *)
   SB_DFF  dff_29_156 (
      .C       (i_clk         ),
      .D       (p2_dl[156]    ),
      .Q       (p3_dl[156]    )
   );
   (* BEL="X2/Y20/lc5" *)
   SB_DFF  dff_2_157 (
      .C       (i_clk         ),
      .D       (p0_dl[158]  ),
      .Q       (p1_dl[157]    )
   );

   (* BEL="X3/Y20/lc5" *)
   SB_DFF  dff_3_157 (
      .C       (i_clk         ),
      .D       (p1_dl[157]    ),
      .Q       (p2_dl[157]    )
   );


   (* BEL="X29/Y20/lc5" *)
   SB_DFF  dff_29_157 (
      .C       (i_clk         ),
      .D       (p2_dl[157]    ),
      .Q       (p3_dl[157]    )
   );
   (* BEL="X2/Y20/lc6" *)
   SB_DFF  dff_2_158 (
      .C       (i_clk         ),
      .D       (p0_dl[159]  ),
      .Q       (p1_dl[158]    )
   );

   (* BEL="X3/Y20/lc6" *)
   SB_DFF  dff_3_158 (
      .C       (i_clk         ),
      .D       (p1_dl[158]    ),
      .Q       (p2_dl[158]    )
   );


   (* BEL="X29/Y20/lc6" *)
   SB_DFF  dff_29_158 (
      .C       (i_clk         ),
      .D       (p2_dl[158]    ),
      .Q       (p3_dl[158]    )
   );
   (* BEL="X2/Y20/lc7" *)
   SB_DFF  dff_2_159 (
      .C       (i_clk         ),
      .D       (p0_dl[160]  ),
      .Q       (p1_dl[159]    )
   );

   (* BEL="X3/Y20/lc7" *)
   SB_DFF  dff_3_159 (
      .C       (i_clk         ),
      .D       (p1_dl[159]    ),
      .Q       (p2_dl[159]    )
   );


   (* BEL="X29/Y20/lc7" *)
   SB_DFF  dff_29_159 (
      .C       (i_clk         ),
      .D       (p2_dl[159]    ),
      .Q       (p3_dl[159]    )
   );
   (* BEL="X2/Y21/lc0" *)
   SB_DFF  dff_2_160 (
      .C       (i_clk         ),
      .D       (p0_dl[161]  ),
      .Q       (p1_dl[160]    )
   );

   (* BEL="X3/Y21/lc0" *)
   SB_DFF  dff_3_160 (
      .C       (i_clk         ),
      .D       (p1_dl[160]    ),
      .Q       (p2_dl[160]    )
   );


   (* BEL="X29/Y21/lc0" *)
   SB_DFF  dff_29_160 (
      .C       (i_clk         ),
      .D       (p2_dl[160]    ),
      .Q       (p3_dl[160]    )
   );
   (* BEL="X2/Y21/lc1" *)
   SB_DFF  dff_2_161 (
      .C       (i_clk         ),
      .D       (p0_dl[162]  ),
      .Q       (p1_dl[161]    )
   );

   (* BEL="X3/Y21/lc1" *)
   SB_DFF  dff_3_161 (
      .C       (i_clk         ),
      .D       (p1_dl[161]    ),
      .Q       (p2_dl[161]    )
   );


   (* BEL="X29/Y21/lc1" *)
   SB_DFF  dff_29_161 (
      .C       (i_clk         ),
      .D       (p2_dl[161]    ),
      .Q       (p3_dl[161]    )
   );
   (* BEL="X2/Y21/lc2" *)
   SB_DFF  dff_2_162 (
      .C       (i_clk         ),
      .D       (p0_dl[163]  ),
      .Q       (p1_dl[162]    )
   );

   (* BEL="X3/Y21/lc2" *)
   SB_DFF  dff_3_162 (
      .C       (i_clk         ),
      .D       (p1_dl[162]    ),
      .Q       (p2_dl[162]    )
   );


   (* BEL="X29/Y21/lc2" *)
   SB_DFF  dff_29_162 (
      .C       (i_clk         ),
      .D       (p2_dl[162]    ),
      .Q       (p3_dl[162]    )
   );
   (* BEL="X2/Y21/lc3" *)
   SB_DFF  dff_2_163 (
      .C       (i_clk         ),
      .D       (p0_dl[164]  ),
      .Q       (p1_dl[163]    )
   );

   (* BEL="X3/Y21/lc3" *)
   SB_DFF  dff_3_163 (
      .C       (i_clk         ),
      .D       (p1_dl[163]    ),
      .Q       (p2_dl[163]    )
   );


   (* BEL="X29/Y21/lc3" *)
   SB_DFF  dff_29_163 (
      .C       (i_clk         ),
      .D       (p2_dl[163]    ),
      .Q       (p3_dl[163]    )
   );
   (* BEL="X2/Y21/lc4" *)
   SB_DFF  dff_2_164 (
      .C       (i_clk         ),
      .D       (p0_dl[165]  ),
      .Q       (p1_dl[164]    )
   );

   (* BEL="X3/Y21/lc4" *)
   SB_DFF  dff_3_164 (
      .C       (i_clk         ),
      .D       (p1_dl[164]    ),
      .Q       (p2_dl[164]    )
   );


   (* BEL="X29/Y21/lc4" *)
   SB_DFF  dff_29_164 (
      .C       (i_clk         ),
      .D       (p2_dl[164]    ),
      .Q       (p3_dl[164]    )
   );
   (* BEL="X2/Y21/lc5" *)
   SB_DFF  dff_2_165 (
      .C       (i_clk         ),
      .D       (p0_dl[166]  ),
      .Q       (p1_dl[165]    )
   );

   (* BEL="X3/Y21/lc5" *)
   SB_DFF  dff_3_165 (
      .C       (i_clk         ),
      .D       (p1_dl[165]    ),
      .Q       (p2_dl[165]    )
   );


   (* BEL="X29/Y21/lc5" *)
   SB_DFF  dff_29_165 (
      .C       (i_clk         ),
      .D       (p2_dl[165]    ),
      .Q       (p3_dl[165]    )
   );
   (* BEL="X2/Y21/lc6" *)
   SB_DFF  dff_2_166 (
      .C       (i_clk         ),
      .D       (p0_dl[167]  ),
      .Q       (p1_dl[166]    )
   );

   (* BEL="X3/Y21/lc6" *)
   SB_DFF  dff_3_166 (
      .C       (i_clk         ),
      .D       (p1_dl[166]    ),
      .Q       (p2_dl[166]    )
   );


   (* BEL="X29/Y21/lc6" *)
   SB_DFF  dff_29_166 (
      .C       (i_clk         ),
      .D       (p2_dl[166]    ),
      .Q       (p3_dl[166]    )
   );
   (* BEL="X2/Y21/lc7" *)
   SB_DFF  dff_2_167 (
      .C       (i_clk         ),
      .D       (p0_dl[168]  ),
      .Q       (p1_dl[167]    )
   );

   (* BEL="X3/Y21/lc7" *)
   SB_DFF  dff_3_167 (
      .C       (i_clk         ),
      .D       (p1_dl[167]    ),
      .Q       (p2_dl[167]    )
   );


   (* BEL="X29/Y21/lc7" *)
   SB_DFF  dff_29_167 (
      .C       (i_clk         ),
      .D       (p2_dl[167]    ),
      .Q       (p3_dl[167]    )
   );
   (* BEL="X2/Y22/lc0" *)
   SB_DFF  dff_2_168 (
      .C       (i_clk         ),
      .D       (p0_dl[169]  ),
      .Q       (p1_dl[168]    )
   );

   (* BEL="X3/Y22/lc0" *)
   SB_DFF  dff_3_168 (
      .C       (i_clk         ),
      .D       (p1_dl[168]    ),
      .Q       (p2_dl[168]    )
   );


   (* BEL="X29/Y22/lc0" *)
   SB_DFF  dff_29_168 (
      .C       (i_clk         ),
      .D       (p2_dl[168]    ),
      .Q       (p3_dl[168]    )
   );
   (* BEL="X2/Y22/lc1" *)
   SB_DFF  dff_2_169 (
      .C       (i_clk         ),
      .D       (p0_dl[170]  ),
      .Q       (p1_dl[169]    )
   );

   (* BEL="X3/Y22/lc1" *)
   SB_DFF  dff_3_169 (
      .C       (i_clk         ),
      .D       (p1_dl[169]    ),
      .Q       (p2_dl[169]    )
   );


   (* BEL="X29/Y22/lc1" *)
   SB_DFF  dff_29_169 (
      .C       (i_clk         ),
      .D       (p2_dl[169]    ),
      .Q       (p3_dl[169]    )
   );
   (* BEL="X2/Y22/lc2" *)
   SB_DFF  dff_2_170 (
      .C       (i_clk         ),
      .D       (p0_dl[171]  ),
      .Q       (p1_dl[170]    )
   );

   (* BEL="X3/Y22/lc2" *)
   SB_DFF  dff_3_170 (
      .C       (i_clk         ),
      .D       (p1_dl[170]    ),
      .Q       (p2_dl[170]    )
   );


   (* BEL="X29/Y22/lc2" *)
   SB_DFF  dff_29_170 (
      .C       (i_clk         ),
      .D       (p2_dl[170]    ),
      .Q       (p3_dl[170]    )
   );
   (* BEL="X2/Y22/lc3" *)
   SB_DFF  dff_2_171 (
      .C       (i_clk         ),
      .D       (p0_dl[172]  ),
      .Q       (p1_dl[171]    )
   );

   (* BEL="X3/Y22/lc3" *)
   SB_DFF  dff_3_171 (
      .C       (i_clk         ),
      .D       (p1_dl[171]    ),
      .Q       (p2_dl[171]    )
   );


   (* BEL="X29/Y22/lc3" *)
   SB_DFF  dff_29_171 (
      .C       (i_clk         ),
      .D       (p2_dl[171]    ),
      .Q       (p3_dl[171]    )
   );
   (* BEL="X2/Y22/lc4" *)
   SB_DFF  dff_2_172 (
      .C       (i_clk         ),
      .D       (p0_dl[173]  ),
      .Q       (p1_dl[172]    )
   );

   (* BEL="X3/Y22/lc4" *)
   SB_DFF  dff_3_172 (
      .C       (i_clk         ),
      .D       (p1_dl[172]    ),
      .Q       (p2_dl[172]    )
   );


   (* BEL="X29/Y22/lc4" *)
   SB_DFF  dff_29_172 (
      .C       (i_clk         ),
      .D       (p2_dl[172]    ),
      .Q       (p3_dl[172]    )
   );
   (* BEL="X2/Y22/lc5" *)
   SB_DFF  dff_2_173 (
      .C       (i_clk         ),
      .D       (p0_dl[174]  ),
      .Q       (p1_dl[173]    )
   );

   (* BEL="X3/Y22/lc5" *)
   SB_DFF  dff_3_173 (
      .C       (i_clk         ),
      .D       (p1_dl[173]    ),
      .Q       (p2_dl[173]    )
   );


   (* BEL="X29/Y22/lc5" *)
   SB_DFF  dff_29_173 (
      .C       (i_clk         ),
      .D       (p2_dl[173]    ),
      .Q       (p3_dl[173]    )
   );
   (* BEL="X2/Y22/lc6" *)
   SB_DFF  dff_2_174 (
      .C       (i_clk         ),
      .D       (p0_dl[175]  ),
      .Q       (p1_dl[174]    )
   );

   (* BEL="X3/Y22/lc6" *)
   SB_DFF  dff_3_174 (
      .C       (i_clk         ),
      .D       (p1_dl[174]    ),
      .Q       (p2_dl[174]    )
   );


   (* BEL="X29/Y22/lc6" *)
   SB_DFF  dff_29_174 (
      .C       (i_clk         ),
      .D       (p2_dl[174]    ),
      .Q       (p3_dl[174]    )
   );
   (* BEL="X2/Y22/lc7" *)
   SB_DFF  dff_2_175 (
      .C       (i_clk         ),
      .D       (p0_dl[176]  ),
      .Q       (p1_dl[175]    )
   );

   (* BEL="X3/Y22/lc7" *)
   SB_DFF  dff_3_175 (
      .C       (i_clk         ),
      .D       (p1_dl[175]    ),
      .Q       (p2_dl[175]    )
   );


   (* BEL="X29/Y22/lc7" *)
   SB_DFF  dff_29_175 (
      .C       (i_clk         ),
      .D       (p2_dl[175]    ),
      .Q       (p3_dl[175]    )
   );
   (* BEL="X2/Y23/lc0" *)
   SB_DFF  dff_2_176 (
      .C       (i_clk         ),
      .D       (p0_dl[177]  ),
      .Q       (p1_dl[176]    )
   );

   (* BEL="X3/Y23/lc0" *)
   SB_DFF  dff_3_176 (
      .C       (i_clk         ),
      .D       (p1_dl[176]    ),
      .Q       (p2_dl[176]    )
   );


   (* BEL="X29/Y23/lc0" *)
   SB_DFF  dff_29_176 (
      .C       (i_clk         ),
      .D       (p2_dl[176]    ),
      .Q       (p3_dl[176]    )
   );
   (* BEL="X2/Y23/lc1" *)
   SB_DFF  dff_2_177 (
      .C       (i_clk         ),
      .D       (p0_dl[178]  ),
      .Q       (p1_dl[177]    )
   );

   (* BEL="X3/Y23/lc1" *)
   SB_DFF  dff_3_177 (
      .C       (i_clk         ),
      .D       (p1_dl[177]    ),
      .Q       (p2_dl[177]    )
   );


   (* BEL="X29/Y23/lc1" *)
   SB_DFF  dff_29_177 (
      .C       (i_clk         ),
      .D       (p2_dl[177]    ),
      .Q       (p3_dl[177]    )
   );
   (* BEL="X2/Y23/lc2" *)
   SB_DFF  dff_2_178 (
      .C       (i_clk         ),
      .D       (p0_dl[179]  ),
      .Q       (p1_dl[178]    )
   );

   (* BEL="X3/Y23/lc2" *)
   SB_DFF  dff_3_178 (
      .C       (i_clk         ),
      .D       (p1_dl[178]    ),
      .Q       (p2_dl[178]    )
   );


   (* BEL="X29/Y23/lc2" *)
   SB_DFF  dff_29_178 (
      .C       (i_clk         ),
      .D       (p2_dl[178]    ),
      .Q       (p3_dl[178]    )
   );
   (* BEL="X2/Y23/lc3" *)
   SB_DFF  dff_2_179 (
      .C       (i_clk         ),
      .D       (p0_dl[180]  ),
      .Q       (p1_dl[179]    )
   );

   (* BEL="X3/Y23/lc3" *)
   SB_DFF  dff_3_179 (
      .C       (i_clk         ),
      .D       (p1_dl[179]    ),
      .Q       (p2_dl[179]    )
   );


   (* BEL="X29/Y23/lc3" *)
   SB_DFF  dff_29_179 (
      .C       (i_clk         ),
      .D       (p2_dl[179]    ),
      .Q       (p3_dl[179]    )
   );
   (* BEL="X2/Y23/lc4" *)
   SB_DFF  dff_2_180 (
      .C       (i_clk         ),
      .D       (p0_dl[181]  ),
      .Q       (p1_dl[180]    )
   );

   (* BEL="X3/Y23/lc4" *)
   SB_DFF  dff_3_180 (
      .C       (i_clk         ),
      .D       (p1_dl[180]    ),
      .Q       (p2_dl[180]    )
   );


   (* BEL="X29/Y23/lc4" *)
   SB_DFF  dff_29_180 (
      .C       (i_clk         ),
      .D       (p2_dl[180]    ),
      .Q       (p3_dl[180]    )
   );
   (* BEL="X2/Y23/lc5" *)
   SB_DFF  dff_2_181 (
      .C       (i_clk         ),
      .D       (p0_dl[182]  ),
      .Q       (p1_dl[181]    )
   );

   (* BEL="X3/Y23/lc5" *)
   SB_DFF  dff_3_181 (
      .C       (i_clk         ),
      .D       (p1_dl[181]    ),
      .Q       (p2_dl[181]    )
   );


   (* BEL="X29/Y23/lc5" *)
   SB_DFF  dff_29_181 (
      .C       (i_clk         ),
      .D       (p2_dl[181]    ),
      .Q       (p3_dl[181]    )
   );
   (* BEL="X2/Y23/lc6" *)
   SB_DFF  dff_2_182 (
      .C       (i_clk         ),
      .D       (p0_dl[183]  ),
      .Q       (p1_dl[182]    )
   );

   (* BEL="X3/Y23/lc6" *)
   SB_DFF  dff_3_182 (
      .C       (i_clk         ),
      .D       (p1_dl[182]    ),
      .Q       (p2_dl[182]    )
   );


   (* BEL="X29/Y23/lc6" *)
   SB_DFF  dff_29_182 (
      .C       (i_clk         ),
      .D       (p2_dl[182]    ),
      .Q       (p3_dl[182]    )
   );
   (* BEL="X2/Y23/lc7" *)
   SB_DFF  dff_2_183 (
      .C       (i_clk         ),
      .D       (p0_dl[184]  ),
      .Q       (p1_dl[183]    )
   );

   (* BEL="X3/Y23/lc7" *)
   SB_DFF  dff_3_183 (
      .C       (i_clk         ),
      .D       (p1_dl[183]    ),
      .Q       (p2_dl[183]    )
   );


   (* BEL="X29/Y23/lc7" *)
   SB_DFF  dff_29_183 (
      .C       (i_clk         ),
      .D       (p2_dl[183]    ),
      .Q       (p3_dl[183]    )
   );
   (* BEL="X2/Y24/lc0" *)
   SB_DFF  dff_2_184 (
      .C       (i_clk         ),
      .D       (p0_dl[185]  ),
      .Q       (p1_dl[184]    )
   );

   (* BEL="X3/Y24/lc0" *)
   SB_DFF  dff_3_184 (
      .C       (i_clk         ),
      .D       (p1_dl[184]    ),
      .Q       (p2_dl[184]    )
   );


   (* BEL="X29/Y24/lc0" *)
   SB_DFF  dff_29_184 (
      .C       (i_clk         ),
      .D       (p2_dl[184]    ),
      .Q       (p3_dl[184]    )
   );
   (* BEL="X2/Y24/lc1" *)
   SB_DFF  dff_2_185 (
      .C       (i_clk         ),
      .D       (p0_dl[186]  ),
      .Q       (p1_dl[185]    )
   );

   (* BEL="X3/Y24/lc1" *)
   SB_DFF  dff_3_185 (
      .C       (i_clk         ),
      .D       (p1_dl[185]    ),
      .Q       (p2_dl[185]    )
   );


   (* BEL="X29/Y24/lc1" *)
   SB_DFF  dff_29_185 (
      .C       (i_clk         ),
      .D       (p2_dl[185]    ),
      .Q       (p3_dl[185]    )
   );
   (* BEL="X2/Y24/lc2" *)
   SB_DFF  dff_2_186 (
      .C       (i_clk         ),
      .D       (p0_dl[187]  ),
      .Q       (p1_dl[186]    )
   );

   (* BEL="X3/Y24/lc2" *)
   SB_DFF  dff_3_186 (
      .C       (i_clk         ),
      .D       (p1_dl[186]    ),
      .Q       (p2_dl[186]    )
   );


   (* BEL="X29/Y24/lc2" *)
   SB_DFF  dff_29_186 (
      .C       (i_clk         ),
      .D       (p2_dl[186]    ),
      .Q       (p3_dl[186]    )
   );
   (* BEL="X2/Y24/lc3" *)
   SB_DFF  dff_2_187 (
      .C       (i_clk         ),
      .D       (p0_dl[188]  ),
      .Q       (p1_dl[187]    )
   );

   (* BEL="X3/Y24/lc3" *)
   SB_DFF  dff_3_187 (
      .C       (i_clk         ),
      .D       (p1_dl[187]    ),
      .Q       (p2_dl[187]    )
   );


   (* BEL="X29/Y24/lc3" *)
   SB_DFF  dff_29_187 (
      .C       (i_clk         ),
      .D       (p2_dl[187]    ),
      .Q       (p3_dl[187]    )
   );
   (* BEL="X2/Y24/lc4" *)
   SB_DFF  dff_2_188 (
      .C       (i_clk         ),
      .D       (p0_dl[189]  ),
      .Q       (p1_dl[188]    )
   );

   (* BEL="X3/Y24/lc4" *)
   SB_DFF  dff_3_188 (
      .C       (i_clk         ),
      .D       (p1_dl[188]    ),
      .Q       (p2_dl[188]    )
   );


   (* BEL="X29/Y24/lc4" *)
   SB_DFF  dff_29_188 (
      .C       (i_clk         ),
      .D       (p2_dl[188]    ),
      .Q       (p3_dl[188]    )
   );
   (* BEL="X2/Y24/lc5" *)
   SB_DFF  dff_2_189 (
      .C       (i_clk         ),
      .D       (p0_dl[190]  ),
      .Q       (p1_dl[189]    )
   );

   (* BEL="X3/Y24/lc5" *)
   SB_DFF  dff_3_189 (
      .C       (i_clk         ),
      .D       (p1_dl[189]    ),
      .Q       (p2_dl[189]    )
   );


   (* BEL="X29/Y24/lc5" *)
   SB_DFF  dff_29_189 (
      .C       (i_clk         ),
      .D       (p2_dl[189]    ),
      .Q       (p3_dl[189]    )
   );
   (* BEL="X2/Y24/lc6" *)
   SB_DFF  dff_2_190 (
      .C       (i_clk         ),
      .D       (p0_dl[191]  ),
      .Q       (p1_dl[190]    )
   );

   (* BEL="X3/Y24/lc6" *)
   SB_DFF  dff_3_190 (
      .C       (i_clk         ),
      .D       (p1_dl[190]    ),
      .Q       (p2_dl[190]    )
   );


   (* BEL="X29/Y24/lc6" *)
   SB_DFF  dff_29_190 (
      .C       (i_clk         ),
      .D       (p2_dl[190]    ),
      .Q       (p3_dl[190]    )
   );
   (* BEL="X2/Y24/lc7" *)
   SB_DFF  dff_2_191 (
      .C       (i_clk         ),
      .D       (p0_dl[192]  ),
      .Q       (p1_dl[191]    )
   );

   (* BEL="X3/Y24/lc7" *)
   SB_DFF  dff_3_191 (
      .C       (i_clk         ),
      .D       (p1_dl[191]    ),
      .Q       (p2_dl[191]    )
   );


   (* BEL="X29/Y24/lc7" *)
   SB_DFF  dff_29_191 (
      .C       (i_clk         ),
      .D       (p2_dl[191]    ),
      .Q       (p3_dl[191]    )
   );
   (* BEL="X2/Y25/lc0" *)
   SB_DFF  dff_2_192 (
      .C       (i_clk         ),
      .D       (p0_dl[193]  ),
      .Q       (p1_dl[192]    )
   );

   (* BEL="X3/Y25/lc0" *)
   SB_DFF  dff_3_192 (
      .C       (i_clk         ),
      .D       (p1_dl[192]    ),
      .Q       (p2_dl[192]    )
   );


   (* BEL="X29/Y25/lc0" *)
   SB_DFF  dff_29_192 (
      .C       (i_clk         ),
      .D       (p2_dl[192]    ),
      .Q       (p3_dl[192]    )
   );
   (* BEL="X2/Y25/lc1" *)
   SB_DFF  dff_2_193 (
      .C       (i_clk         ),
      .D       (p0_dl[194]  ),
      .Q       (p1_dl[193]    )
   );

   (* BEL="X3/Y25/lc1" *)
   SB_DFF  dff_3_193 (
      .C       (i_clk         ),
      .D       (p1_dl[193]    ),
      .Q       (p2_dl[193]    )
   );


   (* BEL="X29/Y25/lc1" *)
   SB_DFF  dff_29_193 (
      .C       (i_clk         ),
      .D       (p2_dl[193]    ),
      .Q       (p3_dl[193]    )
   );
   (* BEL="X2/Y25/lc2" *)
   SB_DFF  dff_2_194 (
      .C       (i_clk         ),
      .D       (p0_dl[195]  ),
      .Q       (p1_dl[194]    )
   );

   (* BEL="X3/Y25/lc2" *)
   SB_DFF  dff_3_194 (
      .C       (i_clk         ),
      .D       (p1_dl[194]    ),
      .Q       (p2_dl[194]    )
   );


   (* BEL="X29/Y25/lc2" *)
   SB_DFF  dff_29_194 (
      .C       (i_clk         ),
      .D       (p2_dl[194]    ),
      .Q       (p3_dl[194]    )
   );
   (* BEL="X2/Y25/lc3" *)
   SB_DFF  dff_2_195 (
      .C       (i_clk         ),
      .D       (p0_dl[196]  ),
      .Q       (p1_dl[195]    )
   );

   (* BEL="X3/Y25/lc3" *)
   SB_DFF  dff_3_195 (
      .C       (i_clk         ),
      .D       (p1_dl[195]    ),
      .Q       (p2_dl[195]    )
   );


   (* BEL="X29/Y25/lc3" *)
   SB_DFF  dff_29_195 (
      .C       (i_clk         ),
      .D       (p2_dl[195]    ),
      .Q       (p3_dl[195]    )
   );
   (* BEL="X2/Y25/lc4" *)
   SB_DFF  dff_2_196 (
      .C       (i_clk         ),
      .D       (p0_dl[197]  ),
      .Q       (p1_dl[196]    )
   );

   (* BEL="X3/Y25/lc4" *)
   SB_DFF  dff_3_196 (
      .C       (i_clk         ),
      .D       (p1_dl[196]    ),
      .Q       (p2_dl[196]    )
   );


   (* BEL="X29/Y25/lc4" *)
   SB_DFF  dff_29_196 (
      .C       (i_clk         ),
      .D       (p2_dl[196]    ),
      .Q       (p3_dl[196]    )
   );
   (* BEL="X2/Y25/lc5" *)
   SB_DFF  dff_2_197 (
      .C       (i_clk         ),
      .D       (p0_dl[198]  ),
      .Q       (p1_dl[197]    )
   );

   (* BEL="X3/Y25/lc5" *)
   SB_DFF  dff_3_197 (
      .C       (i_clk         ),
      .D       (p1_dl[197]    ),
      .Q       (p2_dl[197]    )
   );


   (* BEL="X29/Y25/lc5" *)
   SB_DFF  dff_29_197 (
      .C       (i_clk         ),
      .D       (p2_dl[197]    ),
      .Q       (p3_dl[197]    )
   );
   (* BEL="X2/Y25/lc6" *)
   SB_DFF  dff_2_198 (
      .C       (i_clk         ),
      .D       (p0_dl[199]  ),
      .Q       (p1_dl[198]    )
   );

   (* BEL="X3/Y25/lc6" *)
   SB_DFF  dff_3_198 (
      .C       (i_clk         ),
      .D       (p1_dl[198]    ),
      .Q       (p2_dl[198]    )
   );


   (* BEL="X29/Y25/lc6" *)
   SB_DFF  dff_29_198 (
      .C       (i_clk         ),
      .D       (p2_dl[198]    ),
      .Q       (p3_dl[198]    )
   );
   (* BEL="X2/Y25/lc7" *)
   SB_DFF  dff_2_199 (
      .C       (i_clk         ),
      .D       (p0_dl[200]  ),
      .Q       (p1_dl[199]    )
   );

   (* BEL="X3/Y25/lc7" *)
   SB_DFF  dff_3_199 (
      .C       (i_clk         ),
      .D       (p1_dl[199]    ),
      .Q       (p2_dl[199]    )
   );


   (* BEL="X29/Y25/lc7" *)
   SB_DFF  dff_29_199 (
      .C       (i_clk         ),
      .D       (p2_dl[199]    ),
      .Q       (p3_dl[199]    )
   );
   (* BEL="X2/Y26/lc0" *)
   SB_DFF  dff_2_200 (
      .C       (i_clk         ),
      .D       (p0_dl[201]  ),
      .Q       (p1_dl[200]    )
   );

   (* BEL="X3/Y26/lc0" *)
   SB_DFF  dff_3_200 (
      .C       (i_clk         ),
      .D       (p1_dl[200]    ),
      .Q       (p2_dl[200]    )
   );


   (* BEL="X29/Y26/lc0" *)
   SB_DFF  dff_29_200 (
      .C       (i_clk         ),
      .D       (p2_dl[200]    ),
      .Q       (p3_dl[200]    )
   );
   (* BEL="X2/Y26/lc1" *)
   SB_DFF  dff_2_201 (
      .C       (i_clk         ),
      .D       (p0_dl[202]  ),
      .Q       (p1_dl[201]    )
   );

   (* BEL="X3/Y26/lc1" *)
   SB_DFF  dff_3_201 (
      .C       (i_clk         ),
      .D       (p1_dl[201]    ),
      .Q       (p2_dl[201]    )
   );


   (* BEL="X29/Y26/lc1" *)
   SB_DFF  dff_29_201 (
      .C       (i_clk         ),
      .D       (p2_dl[201]    ),
      .Q       (p3_dl[201]    )
   );
   (* BEL="X2/Y26/lc2" *)
   SB_DFF  dff_2_202 (
      .C       (i_clk         ),
      .D       (p0_dl[203]  ),
      .Q       (p1_dl[202]    )
   );

   (* BEL="X3/Y26/lc2" *)
   SB_DFF  dff_3_202 (
      .C       (i_clk         ),
      .D       (p1_dl[202]    ),
      .Q       (p2_dl[202]    )
   );


   (* BEL="X29/Y26/lc2" *)
   SB_DFF  dff_29_202 (
      .C       (i_clk         ),
      .D       (p2_dl[202]    ),
      .Q       (p3_dl[202]    )
   );
   (* BEL="X2/Y26/lc3" *)
   SB_DFF  dff_2_203 (
      .C       (i_clk         ),
      .D       (p0_dl[204]  ),
      .Q       (p1_dl[203]    )
   );

   (* BEL="X3/Y26/lc3" *)
   SB_DFF  dff_3_203 (
      .C       (i_clk         ),
      .D       (p1_dl[203]    ),
      .Q       (p2_dl[203]    )
   );


   (* BEL="X29/Y26/lc3" *)
   SB_DFF  dff_29_203 (
      .C       (i_clk         ),
      .D       (p2_dl[203]    ),
      .Q       (p3_dl[203]    )
   );
   (* BEL="X2/Y26/lc4" *)
   SB_DFF  dff_2_204 (
      .C       (i_clk         ),
      .D       (p0_dl[205]  ),
      .Q       (p1_dl[204]    )
   );

   (* BEL="X3/Y26/lc4" *)
   SB_DFF  dff_3_204 (
      .C       (i_clk         ),
      .D       (p1_dl[204]    ),
      .Q       (p2_dl[204]    )
   );


   (* BEL="X29/Y26/lc4" *)
   SB_DFF  dff_29_204 (
      .C       (i_clk         ),
      .D       (p2_dl[204]    ),
      .Q       (p3_dl[204]    )
   );
   (* BEL="X2/Y26/lc5" *)
   SB_DFF  dff_2_205 (
      .C       (i_clk         ),
      .D       (p0_dl[206]  ),
      .Q       (p1_dl[205]    )
   );

   (* BEL="X3/Y26/lc5" *)
   SB_DFF  dff_3_205 (
      .C       (i_clk         ),
      .D       (p1_dl[205]    ),
      .Q       (p2_dl[205]    )
   );


   (* BEL="X29/Y26/lc5" *)
   SB_DFF  dff_29_205 (
      .C       (i_clk         ),
      .D       (p2_dl[205]    ),
      .Q       (p3_dl[205]    )
   );
   (* BEL="X2/Y26/lc6" *)
   SB_DFF  dff_2_206 (
      .C       (i_clk         ),
      .D       (p0_dl[207]  ),
      .Q       (p1_dl[206]    )
   );

   (* BEL="X3/Y26/lc6" *)
   SB_DFF  dff_3_206 (
      .C       (i_clk         ),
      .D       (p1_dl[206]    ),
      .Q       (p2_dl[206]    )
   );


   (* BEL="X29/Y26/lc6" *)
   SB_DFF  dff_29_206 (
      .C       (i_clk         ),
      .D       (p2_dl[206]    ),
      .Q       (p3_dl[206]    )
   );
   (* BEL="X2/Y26/lc7" *)
   SB_DFF  dff_2_207 (
      .C       (i_clk         ),
      .D       (p0_dl[208]  ),
      .Q       (p1_dl[207]    )
   );

   (* BEL="X3/Y26/lc7" *)
   SB_DFF  dff_3_207 (
      .C       (i_clk         ),
      .D       (p1_dl[207]    ),
      .Q       (p2_dl[207]    )
   );


   (* BEL="X29/Y26/lc7" *)
   SB_DFF  dff_29_207 (
      .C       (i_clk         ),
      .D       (p2_dl[207]    ),
      .Q       (p3_dl[207]    )
   );
   (* BEL="X2/Y27/lc0" *)
   SB_DFF  dff_2_208 (
      .C       (i_clk         ),
      .D       (p0_dl[209]  ),
      .Q       (p1_dl[208]    )
   );

   (* BEL="X3/Y27/lc0" *)
   SB_DFF  dff_3_208 (
      .C       (i_clk         ),
      .D       (p1_dl[208]    ),
      .Q       (p2_dl[208]    )
   );


   (* BEL="X29/Y27/lc0" *)
   SB_DFF  dff_29_208 (
      .C       (i_clk         ),
      .D       (p2_dl[208]    ),
      .Q       (p3_dl[208]    )
   );
   (* BEL="X2/Y27/lc1" *)
   SB_DFF  dff_2_209 (
      .C       (i_clk         ),
      .D       (p0_dl[210]  ),
      .Q       (p1_dl[209]    )
   );

   (* BEL="X3/Y27/lc1" *)
   SB_DFF  dff_3_209 (
      .C       (i_clk         ),
      .D       (p1_dl[209]    ),
      .Q       (p2_dl[209]    )
   );


   (* BEL="X29/Y27/lc1" *)
   SB_DFF  dff_29_209 (
      .C       (i_clk         ),
      .D       (p2_dl[209]    ),
      .Q       (p3_dl[209]    )
   );
   (* BEL="X2/Y27/lc2" *)
   SB_DFF  dff_2_210 (
      .C       (i_clk         ),
      .D       (p0_dl[211]  ),
      .Q       (p1_dl[210]    )
   );

   (* BEL="X3/Y27/lc2" *)
   SB_DFF  dff_3_210 (
      .C       (i_clk         ),
      .D       (p1_dl[210]    ),
      .Q       (p2_dl[210]    )
   );


   (* BEL="X29/Y27/lc2" *)
   SB_DFF  dff_29_210 (
      .C       (i_clk         ),
      .D       (p2_dl[210]    ),
      .Q       (p3_dl[210]    )
   );
   (* BEL="X2/Y27/lc3" *)
   SB_DFF  dff_2_211 (
      .C       (i_clk         ),
      .D       (p0_dl[212]  ),
      .Q       (p1_dl[211]    )
   );

   (* BEL="X3/Y27/lc3" *)
   SB_DFF  dff_3_211 (
      .C       (i_clk         ),
      .D       (p1_dl[211]    ),
      .Q       (p2_dl[211]    )
   );


   (* BEL="X29/Y27/lc3" *)
   SB_DFF  dff_29_211 (
      .C       (i_clk         ),
      .D       (p2_dl[211]    ),
      .Q       (p3_dl[211]    )
   );
   (* BEL="X2/Y27/lc4" *)
   SB_DFF  dff_2_212 (
      .C       (i_clk         ),
      .D       (p0_dl[213]  ),
      .Q       (p1_dl[212]    )
   );

   (* BEL="X3/Y27/lc4" *)
   SB_DFF  dff_3_212 (
      .C       (i_clk         ),
      .D       (p1_dl[212]    ),
      .Q       (p2_dl[212]    )
   );


   (* BEL="X29/Y27/lc4" *)
   SB_DFF  dff_29_212 (
      .C       (i_clk         ),
      .D       (p2_dl[212]    ),
      .Q       (p3_dl[212]    )
   );
   (* BEL="X2/Y27/lc5" *)
   SB_DFF  dff_2_213 (
      .C       (i_clk         ),
      .D       (p0_dl[214]  ),
      .Q       (p1_dl[213]    )
   );

   (* BEL="X3/Y27/lc5" *)
   SB_DFF  dff_3_213 (
      .C       (i_clk         ),
      .D       (p1_dl[213]    ),
      .Q       (p2_dl[213]    )
   );


   (* BEL="X29/Y27/lc5" *)
   SB_DFF  dff_29_213 (
      .C       (i_clk         ),
      .D       (p2_dl[213]    ),
      .Q       (p3_dl[213]    )
   );
   (* BEL="X2/Y27/lc6" *)
   SB_DFF  dff_2_214 (
      .C       (i_clk         ),
      .D       (p0_dl[215]  ),
      .Q       (p1_dl[214]    )
   );

   (* BEL="X3/Y27/lc6" *)
   SB_DFF  dff_3_214 (
      .C       (i_clk         ),
      .D       (p1_dl[214]    ),
      .Q       (p2_dl[214]    )
   );


   (* BEL="X29/Y27/lc6" *)
   SB_DFF  dff_29_214 (
      .C       (i_clk         ),
      .D       (p2_dl[214]    ),
      .Q       (p3_dl[214]    )
   );
   (* BEL="X2/Y27/lc7" *)
   SB_DFF  dff_2_215 (
      .C       (i_clk         ),
      .D       (p0_dl[216]  ),
      .Q       (p1_dl[215]    )
   );

   (* BEL="X3/Y27/lc7" *)
   SB_DFF  dff_3_215 (
      .C       (i_clk         ),
      .D       (p1_dl[215]    ),
      .Q       (p2_dl[215]    )
   );


   (* BEL="X29/Y27/lc7" *)
   SB_DFF  dff_29_215 (
      .C       (i_clk         ),
      .D       (p2_dl[215]    ),
      .Q       (p3_dl[215]    )
   );
   (* BEL="X2/Y28/lc0" *)
   SB_DFF  dff_2_216 (
      .C       (i_clk         ),
      .D       (p0_dl[217]  ),
      .Q       (p1_dl[216]    )
   );

   (* BEL="X3/Y28/lc0" *)
   SB_DFF  dff_3_216 (
      .C       (i_clk         ),
      .D       (p1_dl[216]    ),
      .Q       (p2_dl[216]    )
   );


   (* BEL="X29/Y28/lc0" *)
   SB_DFF  dff_29_216 (
      .C       (i_clk         ),
      .D       (p2_dl[216]    ),
      .Q       (p3_dl[216]    )
   );
   (* BEL="X2/Y28/lc1" *)
   SB_DFF  dff_2_217 (
      .C       (i_clk         ),
      .D       (p0_dl[218]  ),
      .Q       (p1_dl[217]    )
   );

   (* BEL="X3/Y28/lc1" *)
   SB_DFF  dff_3_217 (
      .C       (i_clk         ),
      .D       (p1_dl[217]    ),
      .Q       (p2_dl[217]    )
   );


   (* BEL="X29/Y28/lc1" *)
   SB_DFF  dff_29_217 (
      .C       (i_clk         ),
      .D       (p2_dl[217]    ),
      .Q       (p3_dl[217]    )
   );
   (* BEL="X2/Y28/lc2" *)
   SB_DFF  dff_2_218 (
      .C       (i_clk         ),
      .D       (p0_dl[219]  ),
      .Q       (p1_dl[218]    )
   );

   (* BEL="X3/Y28/lc2" *)
   SB_DFF  dff_3_218 (
      .C       (i_clk         ),
      .D       (p1_dl[218]    ),
      .Q       (p2_dl[218]    )
   );


   (* BEL="X29/Y28/lc2" *)
   SB_DFF  dff_29_218 (
      .C       (i_clk         ),
      .D       (p2_dl[218]    ),
      .Q       (p3_dl[218]    )
   );
   (* BEL="X2/Y28/lc3" *)
   SB_DFF  dff_2_219 (
      .C       (i_clk         ),
      .D       (p0_dl[220]  ),
      .Q       (p1_dl[219]    )
   );

   (* BEL="X3/Y28/lc3" *)
   SB_DFF  dff_3_219 (
      .C       (i_clk         ),
      .D       (p1_dl[219]    ),
      .Q       (p2_dl[219]    )
   );


   (* BEL="X29/Y28/lc3" *)
   SB_DFF  dff_29_219 (
      .C       (i_clk         ),
      .D       (p2_dl[219]    ),
      .Q       (p3_dl[219]    )
   );
   (* BEL="X2/Y28/lc4" *)
   SB_DFF  dff_2_220 (
      .C       (i_clk         ),
      .D       (p0_dl[221]  ),
      .Q       (p1_dl[220]    )
   );

   (* BEL="X3/Y28/lc4" *)
   SB_DFF  dff_3_220 (
      .C       (i_clk         ),
      .D       (p1_dl[220]    ),
      .Q       (p2_dl[220]    )
   );


   (* BEL="X29/Y28/lc4" *)
   SB_DFF  dff_29_220 (
      .C       (i_clk         ),
      .D       (p2_dl[220]    ),
      .Q       (p3_dl[220]    )
   );
   (* BEL="X2/Y28/lc5" *)
   SB_DFF  dff_2_221 (
      .C       (i_clk         ),
      .D       (p0_dl[222]  ),
      .Q       (p1_dl[221]    )
   );

   (* BEL="X3/Y28/lc5" *)
   SB_DFF  dff_3_221 (
      .C       (i_clk         ),
      .D       (p1_dl[221]    ),
      .Q       (p2_dl[221]    )
   );


   (* BEL="X29/Y28/lc5" *)
   SB_DFF  dff_29_221 (
      .C       (i_clk         ),
      .D       (p2_dl[221]    ),
      .Q       (p3_dl[221]    )
   );
   (* BEL="X2/Y28/lc6" *)
   SB_DFF  dff_2_222 (
      .C       (i_clk         ),
      .D       (p0_dl[223]  ),
      .Q       (p1_dl[222]    )
   );

   (* BEL="X3/Y28/lc6" *)
   SB_DFF  dff_3_222 (
      .C       (i_clk         ),
      .D       (p1_dl[222]    ),
      .Q       (p2_dl[222]    )
   );


   (* BEL="X29/Y28/lc6" *)
   SB_DFF  dff_29_222 (
      .C       (i_clk         ),
      .D       (p2_dl[222]    ),
      .Q       (p3_dl[222]    )
   );
   (* BEL="X2/Y28/lc7" *)
   SB_DFF  dff_2_223 (
      .C       (i_clk         ),
      .D       (p0_dl[224]  ),
      .Q       (p1_dl[223]    )
   );

   (* BEL="X3/Y28/lc7" *)
   SB_DFF  dff_3_223 (
      .C       (i_clk         ),
      .D       (p1_dl[223]    ),
      .Q       (p2_dl[223]    )
   );


   (* BEL="X29/Y28/lc7" *)
   SB_DFF  dff_29_223 (
      .C       (i_clk         ),
      .D       (p2_dl[223]    ),
      .Q       (p3_dl[223]    )
   );
   (* BEL="X2/Y29/lc0" *)
   SB_DFF  dff_2_224 (
      .C       (i_clk         ),
      .D       (p0_dl[225]  ),
      .Q       (p1_dl[224]    )
   );

   (* BEL="X3/Y29/lc0" *)
   SB_DFF  dff_3_224 (
      .C       (i_clk         ),
      .D       (p1_dl[224]    ),
      .Q       (p2_dl[224]    )
   );


   (* BEL="X29/Y29/lc0" *)
   SB_DFF  dff_29_224 (
      .C       (i_clk         ),
      .D       (p2_dl[224]    ),
      .Q       (p3_dl[224]    )
   );
   (* BEL="X2/Y29/lc1" *)
   SB_DFF  dff_2_225 (
      .C       (i_clk         ),
      .D       (p0_dl[226]  ),
      .Q       (p1_dl[225]    )
   );

   (* BEL="X3/Y29/lc1" *)
   SB_DFF  dff_3_225 (
      .C       (i_clk         ),
      .D       (p1_dl[225]    ),
      .Q       (p2_dl[225]    )
   );


   (* BEL="X29/Y29/lc1" *)
   SB_DFF  dff_29_225 (
      .C       (i_clk         ),
      .D       (p2_dl[225]    ),
      .Q       (p3_dl[225]    )
   );
   (* BEL="X2/Y29/lc2" *)
   SB_DFF  dff_2_226 (
      .C       (i_clk         ),
      .D       (p0_dl[227]  ),
      .Q       (p1_dl[226]    )
   );

   (* BEL="X3/Y29/lc2" *)
   SB_DFF  dff_3_226 (
      .C       (i_clk         ),
      .D       (p1_dl[226]    ),
      .Q       (p2_dl[226]    )
   );


   (* BEL="X29/Y29/lc2" *)
   SB_DFF  dff_29_226 (
      .C       (i_clk         ),
      .D       (p2_dl[226]    ),
      .Q       (p3_dl[226]    )
   );
   (* BEL="X2/Y29/lc3" *)
   SB_DFF  dff_2_227 (
      .C       (i_clk         ),
      .D       (p0_dl[228]  ),
      .Q       (p1_dl[227]    )
   );

   (* BEL="X3/Y29/lc3" *)
   SB_DFF  dff_3_227 (
      .C       (i_clk         ),
      .D       (p1_dl[227]    ),
      .Q       (p2_dl[227]    )
   );


   (* BEL="X29/Y29/lc3" *)
   SB_DFF  dff_29_227 (
      .C       (i_clk         ),
      .D       (p2_dl[227]    ),
      .Q       (p3_dl[227]    )
   );
   (* BEL="X2/Y29/lc4" *)
   SB_DFF  dff_2_228 (
      .C       (i_clk         ),
      .D       (p0_dl[229]  ),
      .Q       (p1_dl[228]    )
   );

   (* BEL="X3/Y29/lc4" *)
   SB_DFF  dff_3_228 (
      .C       (i_clk         ),
      .D       (p1_dl[228]    ),
      .Q       (p2_dl[228]    )
   );


   (* BEL="X29/Y29/lc4" *)
   SB_DFF  dff_29_228 (
      .C       (i_clk         ),
      .D       (p2_dl[228]    ),
      .Q       (p3_dl[228]    )
   );
   (* BEL="X2/Y29/lc5" *)
   SB_DFF  dff_2_229 (
      .C       (i_clk         ),
      .D       (p0_dl[230]  ),
      .Q       (p1_dl[229]    )
   );

   (* BEL="X3/Y29/lc5" *)
   SB_DFF  dff_3_229 (
      .C       (i_clk         ),
      .D       (p1_dl[229]    ),
      .Q       (p2_dl[229]    )
   );


   (* BEL="X29/Y29/lc5" *)
   SB_DFF  dff_29_229 (
      .C       (i_clk         ),
      .D       (p2_dl[229]    ),
      .Q       (p3_dl[229]    )
   );
   (* BEL="X2/Y29/lc6" *)
   SB_DFF  dff_2_230 (
      .C       (i_clk         ),
      .D       (p0_dl[231]  ),
      .Q       (p1_dl[230]    )
   );

   (* BEL="X3/Y29/lc6" *)
   SB_DFF  dff_3_230 (
      .C       (i_clk         ),
      .D       (p1_dl[230]    ),
      .Q       (p2_dl[230]    )
   );


   (* BEL="X29/Y29/lc6" *)
   SB_DFF  dff_29_230 (
      .C       (i_clk         ),
      .D       (p2_dl[230]    ),
      .Q       (p3_dl[230]    )
   );
   (* BEL="X2/Y29/lc7" *)
   SB_DFF  dff_2_231 (
      .C       (i_clk         ),
      .D       (p0_dl[232]  ),
      .Q       (p1_dl[231]    )
   );

   (* BEL="X3/Y29/lc7" *)
   SB_DFF  dff_3_231 (
      .C       (i_clk         ),
      .D       (p1_dl[231]    ),
      .Q       (p2_dl[231]    )
   );


   (* BEL="X29/Y29/lc7" *)
   SB_DFF  dff_29_231 (
      .C       (i_clk         ),
      .D       (p2_dl[231]    ),
      .Q       (p3_dl[231]    )
   );
   (* BEL="X2/Y30/lc0" *)
   SB_DFF  dff_2_232 (
      .C       (i_clk         ),
      .D       (p0_dl[233]  ),
      .Q       (p1_dl[232]    )
   );

   (* BEL="X3/Y30/lc0" *)
   SB_DFF  dff_3_232 (
      .C       (i_clk         ),
      .D       (p1_dl[232]    ),
      .Q       (p2_dl[232]    )
   );


   (* BEL="X29/Y30/lc0" *)
   SB_DFF  dff_29_232 (
      .C       (i_clk         ),
      .D       (p2_dl[232]    ),
      .Q       (p3_dl[232]    )
   );
   (* BEL="X2/Y30/lc1" *)
   SB_DFF  dff_2_233 (
      .C       (i_clk         ),
      .D       (p0_dl[234]  ),
      .Q       (p1_dl[233]    )
   );

   (* BEL="X3/Y30/lc1" *)
   SB_DFF  dff_3_233 (
      .C       (i_clk         ),
      .D       (p1_dl[233]    ),
      .Q       (p2_dl[233]    )
   );


   (* BEL="X29/Y30/lc1" *)
   SB_DFF  dff_29_233 (
      .C       (i_clk         ),
      .D       (p2_dl[233]    ),
      .Q       (p3_dl[233]    )
   );
   (* BEL="X2/Y30/lc2" *)
   SB_DFF  dff_2_234 (
      .C       (i_clk         ),
      .D       (p0_dl[235]  ),
      .Q       (p1_dl[234]    )
   );

   (* BEL="X3/Y30/lc2" *)
   SB_DFF  dff_3_234 (
      .C       (i_clk         ),
      .D       (p1_dl[234]    ),
      .Q       (p2_dl[234]    )
   );


   (* BEL="X29/Y30/lc2" *)
   SB_DFF  dff_29_234 (
      .C       (i_clk         ),
      .D       (p2_dl[234]    ),
      .Q       (p3_dl[234]    )
   );
   (* BEL="X2/Y30/lc3" *)
   SB_DFF  dff_2_235 (
      .C       (i_clk         ),
      .D       (p0_dl[236]  ),
      .Q       (p1_dl[235]    )
   );

   (* BEL="X3/Y30/lc3" *)
   SB_DFF  dff_3_235 (
      .C       (i_clk         ),
      .D       (p1_dl[235]    ),
      .Q       (p2_dl[235]    )
   );


   (* BEL="X29/Y30/lc3" *)
   SB_DFF  dff_29_235 (
      .C       (i_clk         ),
      .D       (p2_dl[235]    ),
      .Q       (p3_dl[235]    )
   );
   (* BEL="X2/Y30/lc4" *)
   SB_DFF  dff_2_236 (
      .C       (i_clk         ),
      .D       (p0_dl[237]  ),
      .Q       (p1_dl[236]    )
   );

   (* BEL="X3/Y30/lc4" *)
   SB_DFF  dff_3_236 (
      .C       (i_clk         ),
      .D       (p1_dl[236]    ),
      .Q       (p2_dl[236]    )
   );


   (* BEL="X29/Y30/lc4" *)
   SB_DFF  dff_29_236 (
      .C       (i_clk         ),
      .D       (p2_dl[236]    ),
      .Q       (p3_dl[236]    )
   );
   (* BEL="X2/Y30/lc5" *)
   SB_DFF  dff_2_237 (
      .C       (i_clk         ),
      .D       (p0_dl[238]  ),
      .Q       (p1_dl[237]    )
   );

   (* BEL="X3/Y30/lc5" *)
   SB_DFF  dff_3_237 (
      .C       (i_clk         ),
      .D       (p1_dl[237]    ),
      .Q       (p2_dl[237]    )
   );


   (* BEL="X29/Y30/lc5" *)
   SB_DFF  dff_29_237 (
      .C       (i_clk         ),
      .D       (p2_dl[237]    ),
      .Q       (p3_dl[237]    )
   );
   (* BEL="X2/Y30/lc6" *)
   SB_DFF  dff_2_238 (
      .C       (i_clk         ),
      .D       (p0_dl[239]  ),
      .Q       (p1_dl[238]    )
   );

   (* BEL="X3/Y30/lc6" *)
   SB_DFF  dff_3_238 (
      .C       (i_clk         ),
      .D       (p1_dl[238]    ),
      .Q       (p2_dl[238]    )
   );


   (* BEL="X29/Y30/lc6" *)
   SB_DFF  dff_29_238 (
      .C       (i_clk         ),
      .D       (p2_dl[238]    ),
      .Q       (p3_dl[238]    )
   );
   (* BEL="X2/Y30/lc7" *)
   SB_DFF  dff_2_239 (
      .C       (i_clk         ),
      .D       (p0_dl[240]  ),
      .Q       (p1_dl[239]    )
   );

   (* BEL="X3/Y30/lc7" *)
   SB_DFF  dff_3_239 (
      .C       (i_clk         ),
      .D       (p1_dl[239]    ),
      .Q       (p2_dl[239]    )
   );


   (* BEL="X29/Y30/lc7" *)
   SB_DFF  dff_29_239 (
      .C       (i_clk         ),
      .D       (p2_dl[239]    ),
      .Q       (p3_dl[239]    )
   );
   (* BEL="X2/Y31/lc0" *)
   SB_DFF  dff_2_240 (
      .C       (i_clk         ),
      .D       (p0_dl[241]  ),
      .Q       (p1_dl[240]    )
   );

   (* BEL="X3/Y31/lc0" *)
   SB_DFF  dff_3_240 (
      .C       (i_clk         ),
      .D       (p1_dl[240]    ),
      .Q       (p2_dl[240]    )
   );


   (* BEL="X29/Y31/lc0" *)
   SB_DFF  dff_29_240 (
      .C       (i_clk         ),
      .D       (p2_dl[240]    ),
      .Q       (p3_dl[240]    )
   );
   (* BEL="X2/Y31/lc1" *)
   SB_DFF  dff_2_241 (
      .C       (i_clk         ),
      .D       (p0_dl[242]  ),
      .Q       (p1_dl[241]    )
   );

   (* BEL="X3/Y31/lc1" *)
   SB_DFF  dff_3_241 (
      .C       (i_clk         ),
      .D       (p1_dl[241]    ),
      .Q       (p2_dl[241]    )
   );


   (* BEL="X29/Y31/lc1" *)
   SB_DFF  dff_29_241 (
      .C       (i_clk         ),
      .D       (p2_dl[241]    ),
      .Q       (p3_dl[241]    )
   );
   (* BEL="X2/Y31/lc2" *)
   SB_DFF  dff_2_242 (
      .C       (i_clk         ),
      .D       (p0_dl[243]  ),
      .Q       (p1_dl[242]    )
   );

   (* BEL="X3/Y31/lc2" *)
   SB_DFF  dff_3_242 (
      .C       (i_clk         ),
      .D       (p1_dl[242]    ),
      .Q       (p2_dl[242]    )
   );


   (* BEL="X29/Y31/lc2" *)
   SB_DFF  dff_29_242 (
      .C       (i_clk         ),
      .D       (p2_dl[242]    ),
      .Q       (p3_dl[242]    )
   );
   (* BEL="X2/Y31/lc3" *)
   SB_DFF  dff_2_243 (
      .C       (i_clk         ),
      .D       (p0_dl[244]  ),
      .Q       (p1_dl[243]    )
   );

   (* BEL="X3/Y31/lc3" *)
   SB_DFF  dff_3_243 (
      .C       (i_clk         ),
      .D       (p1_dl[243]    ),
      .Q       (p2_dl[243]    )
   );


   (* BEL="X29/Y31/lc3" *)
   SB_DFF  dff_29_243 (
      .C       (i_clk         ),
      .D       (p2_dl[243]    ),
      .Q       (p3_dl[243]    )
   );
   (* BEL="X2/Y31/lc4" *)
   SB_DFF  dff_2_244 (
      .C       (i_clk         ),
      .D       (p0_dl[245]  ),
      .Q       (p1_dl[244]    )
   );

   (* BEL="X3/Y31/lc4" *)
   SB_DFF  dff_3_244 (
      .C       (i_clk         ),
      .D       (p1_dl[244]    ),
      .Q       (p2_dl[244]    )
   );


   (* BEL="X29/Y31/lc4" *)
   SB_DFF  dff_29_244 (
      .C       (i_clk         ),
      .D       (p2_dl[244]    ),
      .Q       (p3_dl[244]    )
   );
   (* BEL="X2/Y31/lc5" *)
   SB_DFF  dff_2_245 (
      .C       (i_clk         ),
      .D       (p0_dl[246]  ),
      .Q       (p1_dl[245]    )
   );

   (* BEL="X3/Y31/lc5" *)
   SB_DFF  dff_3_245 (
      .C       (i_clk         ),
      .D       (p1_dl[245]    ),
      .Q       (p2_dl[245]    )
   );


   (* BEL="X29/Y31/lc5" *)
   SB_DFF  dff_29_245 (
      .C       (i_clk         ),
      .D       (p2_dl[245]    ),
      .Q       (p3_dl[245]    )
   );
   (* BEL="X2/Y31/lc6" *)
   SB_DFF  dff_2_246 (
      .C       (i_clk         ),
      .D       (p0_dl[247]  ),
      .Q       (p1_dl[246]    )
   );

   (* BEL="X3/Y31/lc6" *)
   SB_DFF  dff_3_246 (
      .C       (i_clk         ),
      .D       (p1_dl[246]    ),
      .Q       (p2_dl[246]    )
   );


   (* BEL="X29/Y31/lc6" *)
   SB_DFF  dff_29_246 (
      .C       (i_clk         ),
      .D       (p2_dl[246]    ),
      .Q       (p3_dl[246]    )
   );
   (* BEL="X2/Y31/lc7" *)
   SB_DFF  dff_2_247 (
      .C       (i_clk         ),
      .D       (p0_dl[248]  ),
      .Q       (p1_dl[247]    )
   );

   (* BEL="X3/Y31/lc7" *)
   SB_DFF  dff_3_247 (
      .C       (i_clk         ),
      .D       (p1_dl[247]    ),
      .Q       (p2_dl[247]    )
   );


   (* BEL="X29/Y31/lc7" *)
   SB_DFF  dff_29_247 (
      .C       (i_clk         ),
      .D       (p2_dl[247]    ),
      .Q       (p3_dl[247]    )
   );
   (* BEL="X2/Y32/lc0" *)
   SB_DFF  dff_2_248 (
      .C       (i_clk         ),
      .D       (p0_dl[249]  ),
      .Q       (p1_dl[248]    )
   );

   (* BEL="X3/Y32/lc0" *)
   SB_DFF  dff_3_248 (
      .C       (i_clk         ),
      .D       (p1_dl[248]    ),
      .Q       (p2_dl[248]    )
   );


   (* BEL="X29/Y32/lc0" *)
   SB_DFF  dff_29_248 (
      .C       (i_clk         ),
      .D       (p2_dl[248]    ),
      .Q       (p3_dl[248]    )
   );
   (* BEL="X2/Y32/lc1" *)
   SB_DFF  dff_2_249 (
      .C       (i_clk         ),
      .D       (p0_dl[250]  ),
      .Q       (p1_dl[249]    )
   );

   (* BEL="X3/Y32/lc1" *)
   SB_DFF  dff_3_249 (
      .C       (i_clk         ),
      .D       (p1_dl[249]    ),
      .Q       (p2_dl[249]    )
   );


   (* BEL="X29/Y32/lc1" *)
   SB_DFF  dff_29_249 (
      .C       (i_clk         ),
      .D       (p2_dl[249]    ),
      .Q       (p3_dl[249]    )
   );
   (* BEL="X2/Y32/lc2" *)
   SB_DFF  dff_2_250 (
      .C       (i_clk         ),
      .D       (p0_dl[251]  ),
      .Q       (p1_dl[250]    )
   );

   (* BEL="X3/Y32/lc2" *)
   SB_DFF  dff_3_250 (
      .C       (i_clk         ),
      .D       (p1_dl[250]    ),
      .Q       (p2_dl[250]    )
   );


   (* BEL="X29/Y32/lc2" *)
   SB_DFF  dff_29_250 (
      .C       (i_clk         ),
      .D       (p2_dl[250]    ),
      .Q       (p3_dl[250]    )
   );
   (* BEL="X2/Y32/lc3" *)
   SB_DFF  dff_2_251 (
      .C       (i_clk         ),
      .D       (p0_dl[252]  ),
      .Q       (p1_dl[251]    )
   );

   (* BEL="X3/Y32/lc3" *)
   SB_DFF  dff_3_251 (
      .C       (i_clk         ),
      .D       (p1_dl[251]    ),
      .Q       (p2_dl[251]    )
   );


   (* BEL="X29/Y32/lc3" *)
   SB_DFF  dff_29_251 (
      .C       (i_clk         ),
      .D       (p2_dl[251]    ),
      .Q       (p3_dl[251]    )
   );
   (* BEL="X2/Y32/lc4" *)
   SB_DFF  dff_2_252 (
      .C       (i_clk         ),
      .D       (p0_dl[253]  ),
      .Q       (p1_dl[252]    )
   );

   (* BEL="X3/Y32/lc4" *)
   SB_DFF  dff_3_252 (
      .C       (i_clk         ),
      .D       (p1_dl[252]    ),
      .Q       (p2_dl[252]    )
   );


   (* BEL="X29/Y32/lc4" *)
   SB_DFF  dff_29_252 (
      .C       (i_clk         ),
      .D       (p2_dl[252]    ),
      .Q       (p3_dl[252]    )
   );
   (* BEL="X2/Y32/lc5" *)
   SB_DFF  dff_2_253 (
      .C       (i_clk         ),
      .D       (p0_dl[254]  ),
      .Q       (p1_dl[253]    )
   );

   (* BEL="X3/Y32/lc5" *)
   SB_DFF  dff_3_253 (
      .C       (i_clk         ),
      .D       (p1_dl[253]    ),
      .Q       (p2_dl[253]    )
   );


   (* BEL="X29/Y32/lc5" *)
   SB_DFF  dff_29_253 (
      .C       (i_clk         ),
      .D       (p2_dl[253]    ),
      .Q       (p3_dl[253]    )
   );
   (* BEL="X2/Y32/lc6" *)
   SB_DFF  dff_2_254 (
      .C       (i_clk         ),
      .D       (p0_dl[255]  ),
      .Q       (p1_dl[254]    )
   );

   (* BEL="X3/Y32/lc6" *)
   SB_DFF  dff_3_254 (
      .C       (i_clk         ),
      .D       (p1_dl[254]    ),
      .Q       (p2_dl[254]    )
   );


   (* BEL="X29/Y32/lc6" *)
   SB_DFF  dff_29_254 (
      .C       (i_clk         ),
      .D       (p2_dl[254]    ),
      .Q       (p3_dl[254]    )
   );
   (* BEL="X2/Y32/lc7" *)
   SB_DFF  dff_2_255 (
      .C       (i_clk         ),
      .D       (p0_dl[256]  ),
      .Q       (p1_dl[255]    )
   );

   (* BEL="X3/Y32/lc7" *)
   SB_DFF  dff_3_255 (
      .C       (i_clk         ),
      .D       (p1_dl[255]    ),
      .Q       (p2_dl[255]    )
   );


   (* BEL="X29/Y32/lc7" *)
   SB_DFF  dff_29_255 (
      .C       (i_clk         ),
      .D       (p2_dl[255]    ),
      .Q       (p3_dl[255]    )
   );
assign o_data = p3_dl[i_sel];

endmodule

