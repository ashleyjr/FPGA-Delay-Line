module x_variable_delay_line (
   input    logic                   i_dl,
   input    logic [256-1:0]    i_ctrl,
   output   logic                   o_dl
);

logic [256:0]   out;
logic [256:0]   in;

assign out[0] = i_dl;

   (* BEL="X1/Y1/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut0 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[0]      ),
      .O       (out[1]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y1/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut0 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[1]          ),
      .I1      (in[1]              ),
      .I0      (out[1]             ),
      .O       (in[0]                )
   );
   (* BEL="X1/Y1/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut1 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[1]      ),
      .O       (out[2]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y1/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut1 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[2]          ),
      .I1      (in[2]              ),
      .I0      (out[2]             ),
      .O       (in[1]                )
   );
   (* BEL="X1/Y1/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut2 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[2]      ),
      .O       (out[3]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y1/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut2 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[3]          ),
      .I1      (in[3]              ),
      .I0      (out[3]             ),
      .O       (in[2]                )
   );
   (* BEL="X1/Y1/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut3 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[3]      ),
      .O       (out[4]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y1/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut3 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[4]          ),
      .I1      (in[4]              ),
      .I0      (out[4]             ),
      .O       (in[3]                )
   );
   (* BEL="X1/Y1/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut4 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[4]      ),
      .O       (out[5]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y1/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut4 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[5]          ),
      .I1      (in[5]              ),
      .I0      (out[5]             ),
      .O       (in[4]                )
   );
   (* BEL="X1/Y1/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut5 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[5]      ),
      .O       (out[6]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y1/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut5 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[6]          ),
      .I1      (in[6]              ),
      .I0      (out[6]             ),
      .O       (in[5]                )
   );
   (* BEL="X1/Y1/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut6 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[6]      ),
      .O       (out[7]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y1/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut6 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[7]          ),
      .I1      (in[7]              ),
      .I0      (out[7]             ),
      .O       (in[6]                )
   );
   (* BEL="X1/Y1/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut7 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[7]      ),
      .O       (out[8]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y1/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut7 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[8]          ),
      .I1      (in[8]              ),
      .I0      (out[8]             ),
      .O       (in[7]                )
   );
   (* BEL="X1/Y2/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut8 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[8]      ),
      .O       (out[9]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y2/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut8 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[9]          ),
      .I1      (in[9]              ),
      .I0      (out[9]             ),
      .O       (in[8]                )
   );
   (* BEL="X1/Y2/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut9 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[9]      ),
      .O       (out[10]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y2/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut9 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[10]          ),
      .I1      (in[10]              ),
      .I0      (out[10]             ),
      .O       (in[9]                )
   );
   (* BEL="X1/Y2/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut10 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[10]      ),
      .O       (out[11]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y2/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut10 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[11]          ),
      .I1      (in[11]              ),
      .I0      (out[11]             ),
      .O       (in[10]                )
   );
   (* BEL="X1/Y2/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut11 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[11]      ),
      .O       (out[12]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y2/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut11 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[12]          ),
      .I1      (in[12]              ),
      .I0      (out[12]             ),
      .O       (in[11]                )
   );
   (* BEL="X1/Y2/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut12 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[12]      ),
      .O       (out[13]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y2/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut12 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[13]          ),
      .I1      (in[13]              ),
      .I0      (out[13]             ),
      .O       (in[12]                )
   );
   (* BEL="X1/Y2/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut13 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[13]      ),
      .O       (out[14]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y2/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut13 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[14]          ),
      .I1      (in[14]              ),
      .I0      (out[14]             ),
      .O       (in[13]                )
   );
   (* BEL="X1/Y2/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut14 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[14]      ),
      .O       (out[15]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y2/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut14 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[15]          ),
      .I1      (in[15]              ),
      .I0      (out[15]             ),
      .O       (in[14]                )
   );
   (* BEL="X1/Y2/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut15 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[15]      ),
      .O       (out[16]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y2/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut15 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[16]          ),
      .I1      (in[16]              ),
      .I0      (out[16]             ),
      .O       (in[15]                )
   );
   (* BEL="X1/Y3/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut16 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[16]      ),
      .O       (out[17]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y3/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut16 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[17]          ),
      .I1      (in[17]              ),
      .I0      (out[17]             ),
      .O       (in[16]                )
   );
   (* BEL="X1/Y3/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut17 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[17]      ),
      .O       (out[18]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y3/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut17 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[18]          ),
      .I1      (in[18]              ),
      .I0      (out[18]             ),
      .O       (in[17]                )
   );
   (* BEL="X1/Y3/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut18 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[18]      ),
      .O       (out[19]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y3/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut18 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[19]          ),
      .I1      (in[19]              ),
      .I0      (out[19]             ),
      .O       (in[18]                )
   );
   (* BEL="X1/Y3/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut19 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[19]      ),
      .O       (out[20]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y3/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut19 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[20]          ),
      .I1      (in[20]              ),
      .I0      (out[20]             ),
      .O       (in[19]                )
   );
   (* BEL="X1/Y3/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut20 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[20]      ),
      .O       (out[21]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y3/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut20 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[21]          ),
      .I1      (in[21]              ),
      .I0      (out[21]             ),
      .O       (in[20]                )
   );
   (* BEL="X1/Y3/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut21 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[21]      ),
      .O       (out[22]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y3/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut21 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[22]          ),
      .I1      (in[22]              ),
      .I0      (out[22]             ),
      .O       (in[21]                )
   );
   (* BEL="X1/Y3/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut22 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[22]      ),
      .O       (out[23]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y3/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut22 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[23]          ),
      .I1      (in[23]              ),
      .I0      (out[23]             ),
      .O       (in[22]                )
   );
   (* BEL="X1/Y3/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut23 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[23]      ),
      .O       (out[24]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y3/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut23 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[24]          ),
      .I1      (in[24]              ),
      .I0      (out[24]             ),
      .O       (in[23]                )
   );
   (* BEL="X1/Y4/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut24 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[24]      ),
      .O       (out[25]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y4/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut24 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[25]          ),
      .I1      (in[25]              ),
      .I0      (out[25]             ),
      .O       (in[24]                )
   );
   (* BEL="X1/Y4/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut25 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[25]      ),
      .O       (out[26]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y4/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut25 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[26]          ),
      .I1      (in[26]              ),
      .I0      (out[26]             ),
      .O       (in[25]                )
   );
   (* BEL="X1/Y4/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut26 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[26]      ),
      .O       (out[27]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y4/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut26 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[27]          ),
      .I1      (in[27]              ),
      .I0      (out[27]             ),
      .O       (in[26]                )
   );
   (* BEL="X1/Y4/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut27 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[27]      ),
      .O       (out[28]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y4/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut27 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[28]          ),
      .I1      (in[28]              ),
      .I0      (out[28]             ),
      .O       (in[27]                )
   );
   (* BEL="X1/Y4/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut28 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[28]      ),
      .O       (out[29]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y4/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut28 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[29]          ),
      .I1      (in[29]              ),
      .I0      (out[29]             ),
      .O       (in[28]                )
   );
   (* BEL="X1/Y4/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut29 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[29]      ),
      .O       (out[30]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y4/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut29 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[30]          ),
      .I1      (in[30]              ),
      .I0      (out[30]             ),
      .O       (in[29]                )
   );
   (* BEL="X1/Y4/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut30 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[30]      ),
      .O       (out[31]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y4/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut30 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[31]          ),
      .I1      (in[31]              ),
      .I0      (out[31]             ),
      .O       (in[30]                )
   );
   (* BEL="X1/Y4/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut31 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[31]      ),
      .O       (out[32]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y4/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut31 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[32]          ),
      .I1      (in[32]              ),
      .I0      (out[32]             ),
      .O       (in[31]                )
   );
   (* BEL="X1/Y5/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut32 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[32]      ),
      .O       (out[33]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y5/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut32 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[33]          ),
      .I1      (in[33]              ),
      .I0      (out[33]             ),
      .O       (in[32]                )
   );
   (* BEL="X1/Y5/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut33 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[33]      ),
      .O       (out[34]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y5/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut33 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[34]          ),
      .I1      (in[34]              ),
      .I0      (out[34]             ),
      .O       (in[33]                )
   );
   (* BEL="X1/Y5/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut34 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[34]      ),
      .O       (out[35]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y5/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut34 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[35]          ),
      .I1      (in[35]              ),
      .I0      (out[35]             ),
      .O       (in[34]                )
   );
   (* BEL="X1/Y5/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut35 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[35]      ),
      .O       (out[36]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y5/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut35 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[36]          ),
      .I1      (in[36]              ),
      .I0      (out[36]             ),
      .O       (in[35]                )
   );
   (* BEL="X1/Y5/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut36 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[36]      ),
      .O       (out[37]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y5/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut36 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[37]          ),
      .I1      (in[37]              ),
      .I0      (out[37]             ),
      .O       (in[36]                )
   );
   (* BEL="X1/Y5/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut37 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[37]      ),
      .O       (out[38]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y5/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut37 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[38]          ),
      .I1      (in[38]              ),
      .I0      (out[38]             ),
      .O       (in[37]                )
   );
   (* BEL="X1/Y5/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut38 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[38]      ),
      .O       (out[39]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y5/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut38 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[39]          ),
      .I1      (in[39]              ),
      .I0      (out[39]             ),
      .O       (in[38]                )
   );
   (* BEL="X1/Y5/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut39 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[39]      ),
      .O       (out[40]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y5/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut39 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[40]          ),
      .I1      (in[40]              ),
      .I0      (out[40]             ),
      .O       (in[39]                )
   );
   (* BEL="X1/Y6/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut40 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[40]      ),
      .O       (out[41]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y6/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut40 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[41]          ),
      .I1      (in[41]              ),
      .I0      (out[41]             ),
      .O       (in[40]                )
   );
   (* BEL="X1/Y6/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut41 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[41]      ),
      .O       (out[42]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y6/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut41 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[42]          ),
      .I1      (in[42]              ),
      .I0      (out[42]             ),
      .O       (in[41]                )
   );
   (* BEL="X1/Y6/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut42 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[42]      ),
      .O       (out[43]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y6/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut42 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[43]          ),
      .I1      (in[43]              ),
      .I0      (out[43]             ),
      .O       (in[42]                )
   );
   (* BEL="X1/Y6/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut43 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[43]      ),
      .O       (out[44]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y6/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut43 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[44]          ),
      .I1      (in[44]              ),
      .I0      (out[44]             ),
      .O       (in[43]                )
   );
   (* BEL="X1/Y6/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut44 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[44]      ),
      .O       (out[45]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y6/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut44 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[45]          ),
      .I1      (in[45]              ),
      .I0      (out[45]             ),
      .O       (in[44]                )
   );
   (* BEL="X1/Y6/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut45 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[45]      ),
      .O       (out[46]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y6/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut45 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[46]          ),
      .I1      (in[46]              ),
      .I0      (out[46]             ),
      .O       (in[45]                )
   );
   (* BEL="X1/Y6/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut46 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[46]      ),
      .O       (out[47]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y6/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut46 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[47]          ),
      .I1      (in[47]              ),
      .I0      (out[47]             ),
      .O       (in[46]                )
   );
   (* BEL="X1/Y6/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut47 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[47]      ),
      .O       (out[48]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y6/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut47 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[48]          ),
      .I1      (in[48]              ),
      .I0      (out[48]             ),
      .O       (in[47]                )
   );
   (* BEL="X1/Y7/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut48 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[48]      ),
      .O       (out[49]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y7/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut48 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[49]          ),
      .I1      (in[49]              ),
      .I0      (out[49]             ),
      .O       (in[48]                )
   );
   (* BEL="X1/Y7/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut49 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[49]      ),
      .O       (out[50]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y7/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut49 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[50]          ),
      .I1      (in[50]              ),
      .I0      (out[50]             ),
      .O       (in[49]                )
   );
   (* BEL="X1/Y7/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut50 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[50]      ),
      .O       (out[51]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y7/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut50 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[51]          ),
      .I1      (in[51]              ),
      .I0      (out[51]             ),
      .O       (in[50]                )
   );
   (* BEL="X1/Y7/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut51 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[51]      ),
      .O       (out[52]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y7/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut51 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[52]          ),
      .I1      (in[52]              ),
      .I0      (out[52]             ),
      .O       (in[51]                )
   );
   (* BEL="X1/Y7/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut52 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[52]      ),
      .O       (out[53]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y7/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut52 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[53]          ),
      .I1      (in[53]              ),
      .I0      (out[53]             ),
      .O       (in[52]                )
   );
   (* BEL="X1/Y7/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut53 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[53]      ),
      .O       (out[54]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y7/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut53 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[54]          ),
      .I1      (in[54]              ),
      .I0      (out[54]             ),
      .O       (in[53]                )
   );
   (* BEL="X1/Y7/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut54 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[54]      ),
      .O       (out[55]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y7/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut54 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[55]          ),
      .I1      (in[55]              ),
      .I0      (out[55]             ),
      .O       (in[54]                )
   );
   (* BEL="X1/Y7/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut55 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[55]      ),
      .O       (out[56]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y7/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut55 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[56]          ),
      .I1      (in[56]              ),
      .I0      (out[56]             ),
      .O       (in[55]                )
   );
   (* BEL="X1/Y8/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut56 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[56]      ),
      .O       (out[57]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y8/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut56 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[57]          ),
      .I1      (in[57]              ),
      .I0      (out[57]             ),
      .O       (in[56]                )
   );
   (* BEL="X1/Y8/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut57 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[57]      ),
      .O       (out[58]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y8/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut57 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[58]          ),
      .I1      (in[58]              ),
      .I0      (out[58]             ),
      .O       (in[57]                )
   );
   (* BEL="X1/Y8/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut58 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[58]      ),
      .O       (out[59]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y8/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut58 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[59]          ),
      .I1      (in[59]              ),
      .I0      (out[59]             ),
      .O       (in[58]                )
   );
   (* BEL="X1/Y8/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut59 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[59]      ),
      .O       (out[60]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y8/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut59 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[60]          ),
      .I1      (in[60]              ),
      .I0      (out[60]             ),
      .O       (in[59]                )
   );
   (* BEL="X1/Y8/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut60 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[60]      ),
      .O       (out[61]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y8/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut60 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[61]          ),
      .I1      (in[61]              ),
      .I0      (out[61]             ),
      .O       (in[60]                )
   );
   (* BEL="X1/Y8/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut61 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[61]      ),
      .O       (out[62]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y8/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut61 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[62]          ),
      .I1      (in[62]              ),
      .I0      (out[62]             ),
      .O       (in[61]                )
   );
   (* BEL="X1/Y8/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut62 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[62]      ),
      .O       (out[63]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y8/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut62 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[63]          ),
      .I1      (in[63]              ),
      .I0      (out[63]             ),
      .O       (in[62]                )
   );
   (* BEL="X1/Y8/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut63 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[63]      ),
      .O       (out[64]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y8/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut63 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[64]          ),
      .I1      (in[64]              ),
      .I0      (out[64]             ),
      .O       (in[63]                )
   );
   (* BEL="X1/Y9/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut64 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[64]      ),
      .O       (out[65]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y9/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut64 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[65]          ),
      .I1      (in[65]              ),
      .I0      (out[65]             ),
      .O       (in[64]                )
   );
   (* BEL="X1/Y9/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut65 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[65]      ),
      .O       (out[66]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y9/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut65 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[66]          ),
      .I1      (in[66]              ),
      .I0      (out[66]             ),
      .O       (in[65]                )
   );
   (* BEL="X1/Y9/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut66 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[66]      ),
      .O       (out[67]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y9/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut66 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[67]          ),
      .I1      (in[67]              ),
      .I0      (out[67]             ),
      .O       (in[66]                )
   );
   (* BEL="X1/Y9/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut67 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[67]      ),
      .O       (out[68]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y9/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut67 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[68]          ),
      .I1      (in[68]              ),
      .I0      (out[68]             ),
      .O       (in[67]                )
   );
   (* BEL="X1/Y9/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut68 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[68]      ),
      .O       (out[69]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y9/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut68 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[69]          ),
      .I1      (in[69]              ),
      .I0      (out[69]             ),
      .O       (in[68]                )
   );
   (* BEL="X1/Y9/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut69 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[69]      ),
      .O       (out[70]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y9/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut69 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[70]          ),
      .I1      (in[70]              ),
      .I0      (out[70]             ),
      .O       (in[69]                )
   );
   (* BEL="X1/Y9/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut70 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[70]      ),
      .O       (out[71]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y9/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut70 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[71]          ),
      .I1      (in[71]              ),
      .I0      (out[71]             ),
      .O       (in[70]                )
   );
   (* BEL="X1/Y9/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut71 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[71]      ),
      .O       (out[72]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y9/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut71 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[72]          ),
      .I1      (in[72]              ),
      .I0      (out[72]             ),
      .O       (in[71]                )
   );
   (* BEL="X1/Y10/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut72 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[72]      ),
      .O       (out[73]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y10/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut72 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[73]          ),
      .I1      (in[73]              ),
      .I0      (out[73]             ),
      .O       (in[72]                )
   );
   (* BEL="X1/Y10/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut73 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[73]      ),
      .O       (out[74]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y10/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut73 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[74]          ),
      .I1      (in[74]              ),
      .I0      (out[74]             ),
      .O       (in[73]                )
   );
   (* BEL="X1/Y10/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut74 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[74]      ),
      .O       (out[75]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y10/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut74 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[75]          ),
      .I1      (in[75]              ),
      .I0      (out[75]             ),
      .O       (in[74]                )
   );
   (* BEL="X1/Y10/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut75 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[75]      ),
      .O       (out[76]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y10/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut75 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[76]          ),
      .I1      (in[76]              ),
      .I0      (out[76]             ),
      .O       (in[75]                )
   );
   (* BEL="X1/Y10/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut76 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[76]      ),
      .O       (out[77]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y10/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut76 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[77]          ),
      .I1      (in[77]              ),
      .I0      (out[77]             ),
      .O       (in[76]                )
   );
   (* BEL="X1/Y10/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut77 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[77]      ),
      .O       (out[78]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y10/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut77 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[78]          ),
      .I1      (in[78]              ),
      .I0      (out[78]             ),
      .O       (in[77]                )
   );
   (* BEL="X1/Y10/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut78 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[78]      ),
      .O       (out[79]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y10/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut78 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[79]          ),
      .I1      (in[79]              ),
      .I0      (out[79]             ),
      .O       (in[78]                )
   );
   (* BEL="X1/Y10/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut79 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[79]      ),
      .O       (out[80]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y10/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut79 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[80]          ),
      .I1      (in[80]              ),
      .I0      (out[80]             ),
      .O       (in[79]                )
   );
   (* BEL="X1/Y11/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut80 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[80]      ),
      .O       (out[81]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y11/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut80 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[81]          ),
      .I1      (in[81]              ),
      .I0      (out[81]             ),
      .O       (in[80]                )
   );
   (* BEL="X1/Y11/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut81 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[81]      ),
      .O       (out[82]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y11/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut81 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[82]          ),
      .I1      (in[82]              ),
      .I0      (out[82]             ),
      .O       (in[81]                )
   );
   (* BEL="X1/Y11/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut82 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[82]      ),
      .O       (out[83]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y11/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut82 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[83]          ),
      .I1      (in[83]              ),
      .I0      (out[83]             ),
      .O       (in[82]                )
   );
   (* BEL="X1/Y11/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut83 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[83]      ),
      .O       (out[84]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y11/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut83 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[84]          ),
      .I1      (in[84]              ),
      .I0      (out[84]             ),
      .O       (in[83]                )
   );
   (* BEL="X1/Y11/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut84 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[84]      ),
      .O       (out[85]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y11/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut84 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[85]          ),
      .I1      (in[85]              ),
      .I0      (out[85]             ),
      .O       (in[84]                )
   );
   (* BEL="X1/Y11/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut85 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[85]      ),
      .O       (out[86]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y11/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut85 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[86]          ),
      .I1      (in[86]              ),
      .I0      (out[86]             ),
      .O       (in[85]                )
   );
   (* BEL="X1/Y11/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut86 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[86]      ),
      .O       (out[87]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y11/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut86 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[87]          ),
      .I1      (in[87]              ),
      .I0      (out[87]             ),
      .O       (in[86]                )
   );
   (* BEL="X1/Y11/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut87 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[87]      ),
      .O       (out[88]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y11/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut87 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[88]          ),
      .I1      (in[88]              ),
      .I0      (out[88]             ),
      .O       (in[87]                )
   );
   (* BEL="X1/Y12/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut88 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[88]      ),
      .O       (out[89]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y12/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut88 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[89]          ),
      .I1      (in[89]              ),
      .I0      (out[89]             ),
      .O       (in[88]                )
   );
   (* BEL="X1/Y12/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut89 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[89]      ),
      .O       (out[90]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y12/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut89 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[90]          ),
      .I1      (in[90]              ),
      .I0      (out[90]             ),
      .O       (in[89]                )
   );
   (* BEL="X1/Y12/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut90 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[90]      ),
      .O       (out[91]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y12/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut90 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[91]          ),
      .I1      (in[91]              ),
      .I0      (out[91]             ),
      .O       (in[90]                )
   );
   (* BEL="X1/Y12/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut91 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[91]      ),
      .O       (out[92]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y12/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut91 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[92]          ),
      .I1      (in[92]              ),
      .I0      (out[92]             ),
      .O       (in[91]                )
   );
   (* BEL="X1/Y12/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut92 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[92]      ),
      .O       (out[93]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y12/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut92 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[93]          ),
      .I1      (in[93]              ),
      .I0      (out[93]             ),
      .O       (in[92]                )
   );
   (* BEL="X1/Y12/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut93 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[93]      ),
      .O       (out[94]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y12/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut93 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[94]          ),
      .I1      (in[94]              ),
      .I0      (out[94]             ),
      .O       (in[93]                )
   );
   (* BEL="X1/Y12/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut94 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[94]      ),
      .O       (out[95]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y12/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut94 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[95]          ),
      .I1      (in[95]              ),
      .I0      (out[95]             ),
      .O       (in[94]                )
   );
   (* BEL="X1/Y12/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut95 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[95]      ),
      .O       (out[96]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y12/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut95 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[96]          ),
      .I1      (in[96]              ),
      .I0      (out[96]             ),
      .O       (in[95]                )
   );
   (* BEL="X1/Y13/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut96 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[96]      ),
      .O       (out[97]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y13/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut96 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[97]          ),
      .I1      (in[97]              ),
      .I0      (out[97]             ),
      .O       (in[96]                )
   );
   (* BEL="X1/Y13/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut97 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[97]      ),
      .O       (out[98]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y13/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut97 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[98]          ),
      .I1      (in[98]              ),
      .I0      (out[98]             ),
      .O       (in[97]                )
   );
   (* BEL="X1/Y13/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut98 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[98]      ),
      .O       (out[99]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y13/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut98 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[99]          ),
      .I1      (in[99]              ),
      .I0      (out[99]             ),
      .O       (in[98]                )
   );
   (* BEL="X1/Y13/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut99 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[99]      ),
      .O       (out[100]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y13/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut99 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[100]          ),
      .I1      (in[100]              ),
      .I0      (out[100]             ),
      .O       (in[99]                )
   );
   (* BEL="X1/Y13/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut100 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[100]      ),
      .O       (out[101]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y13/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut100 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[101]          ),
      .I1      (in[101]              ),
      .I0      (out[101]             ),
      .O       (in[100]                )
   );
   (* BEL="X1/Y13/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut101 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[101]      ),
      .O       (out[102]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y13/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut101 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[102]          ),
      .I1      (in[102]              ),
      .I0      (out[102]             ),
      .O       (in[101]                )
   );
   (* BEL="X1/Y13/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut102 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[102]      ),
      .O       (out[103]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y13/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut102 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[103]          ),
      .I1      (in[103]              ),
      .I0      (out[103]             ),
      .O       (in[102]                )
   );
   (* BEL="X1/Y13/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut103 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[103]      ),
      .O       (out[104]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y13/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut103 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[104]          ),
      .I1      (in[104]              ),
      .I0      (out[104]             ),
      .O       (in[103]                )
   );
   (* BEL="X1/Y14/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut104 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[104]      ),
      .O       (out[105]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y14/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut104 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[105]          ),
      .I1      (in[105]              ),
      .I0      (out[105]             ),
      .O       (in[104]                )
   );
   (* BEL="X1/Y14/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut105 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[105]      ),
      .O       (out[106]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y14/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut105 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[106]          ),
      .I1      (in[106]              ),
      .I0      (out[106]             ),
      .O       (in[105]                )
   );
   (* BEL="X1/Y14/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut106 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[106]      ),
      .O       (out[107]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y14/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut106 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[107]          ),
      .I1      (in[107]              ),
      .I0      (out[107]             ),
      .O       (in[106]                )
   );
   (* BEL="X1/Y14/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut107 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[107]      ),
      .O       (out[108]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y14/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut107 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[108]          ),
      .I1      (in[108]              ),
      .I0      (out[108]             ),
      .O       (in[107]                )
   );
   (* BEL="X1/Y14/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut108 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[108]      ),
      .O       (out[109]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y14/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut108 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[109]          ),
      .I1      (in[109]              ),
      .I0      (out[109]             ),
      .O       (in[108]                )
   );
   (* BEL="X1/Y14/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut109 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[109]      ),
      .O       (out[110]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y14/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut109 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[110]          ),
      .I1      (in[110]              ),
      .I0      (out[110]             ),
      .O       (in[109]                )
   );
   (* BEL="X1/Y14/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut110 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[110]      ),
      .O       (out[111]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y14/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut110 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[111]          ),
      .I1      (in[111]              ),
      .I0      (out[111]             ),
      .O       (in[110]                )
   );
   (* BEL="X1/Y14/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut111 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[111]      ),
      .O       (out[112]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y14/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut111 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[112]          ),
      .I1      (in[112]              ),
      .I0      (out[112]             ),
      .O       (in[111]                )
   );
   (* BEL="X1/Y15/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut112 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[112]      ),
      .O       (out[113]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y15/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut112 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[113]          ),
      .I1      (in[113]              ),
      .I0      (out[113]             ),
      .O       (in[112]                )
   );
   (* BEL="X1/Y15/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut113 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[113]      ),
      .O       (out[114]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y15/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut113 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[114]          ),
      .I1      (in[114]              ),
      .I0      (out[114]             ),
      .O       (in[113]                )
   );
   (* BEL="X1/Y15/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut114 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[114]      ),
      .O       (out[115]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y15/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut114 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[115]          ),
      .I1      (in[115]              ),
      .I0      (out[115]             ),
      .O       (in[114]                )
   );
   (* BEL="X1/Y15/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut115 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[115]      ),
      .O       (out[116]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y15/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut115 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[116]          ),
      .I1      (in[116]              ),
      .I0      (out[116]             ),
      .O       (in[115]                )
   );
   (* BEL="X1/Y15/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut116 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[116]      ),
      .O       (out[117]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y15/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut116 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[117]          ),
      .I1      (in[117]              ),
      .I0      (out[117]             ),
      .O       (in[116]                )
   );
   (* BEL="X1/Y15/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut117 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[117]      ),
      .O       (out[118]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y15/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut117 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[118]          ),
      .I1      (in[118]              ),
      .I0      (out[118]             ),
      .O       (in[117]                )
   );
   (* BEL="X1/Y15/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut118 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[118]      ),
      .O       (out[119]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y15/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut118 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[119]          ),
      .I1      (in[119]              ),
      .I0      (out[119]             ),
      .O       (in[118]                )
   );
   (* BEL="X1/Y15/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut119 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[119]      ),
      .O       (out[120]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y15/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut119 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[120]          ),
      .I1      (in[120]              ),
      .I0      (out[120]             ),
      .O       (in[119]                )
   );
   (* BEL="X1/Y16/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut120 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[120]      ),
      .O       (out[121]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y16/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut120 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[121]          ),
      .I1      (in[121]              ),
      .I0      (out[121]             ),
      .O       (in[120]                )
   );
   (* BEL="X1/Y16/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut121 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[121]      ),
      .O       (out[122]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y16/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut121 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[122]          ),
      .I1      (in[122]              ),
      .I0      (out[122]             ),
      .O       (in[121]                )
   );
   (* BEL="X1/Y16/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut122 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[122]      ),
      .O       (out[123]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y16/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut122 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[123]          ),
      .I1      (in[123]              ),
      .I0      (out[123]             ),
      .O       (in[122]                )
   );
   (* BEL="X1/Y16/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut123 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[123]      ),
      .O       (out[124]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y16/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut123 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[124]          ),
      .I1      (in[124]              ),
      .I0      (out[124]             ),
      .O       (in[123]                )
   );
   (* BEL="X1/Y16/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut124 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[124]      ),
      .O       (out[125]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y16/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut124 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[125]          ),
      .I1      (in[125]              ),
      .I0      (out[125]             ),
      .O       (in[124]                )
   );
   (* BEL="X1/Y16/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut125 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[125]      ),
      .O       (out[126]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y16/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut125 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[126]          ),
      .I1      (in[126]              ),
      .I0      (out[126]             ),
      .O       (in[125]                )
   );
   (* BEL="X1/Y16/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut126 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[126]      ),
      .O       (out[127]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y16/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut126 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[127]          ),
      .I1      (in[127]              ),
      .I0      (out[127]             ),
      .O       (in[126]                )
   );
   (* BEL="X1/Y16/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut127 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[127]      ),
      .O       (out[128]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y16/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut127 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[128]          ),
      .I1      (in[128]              ),
      .I0      (out[128]             ),
      .O       (in[127]                )
   );
   (* BEL="X1/Y17/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut128 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[128]      ),
      .O       (out[129]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y17/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut128 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[129]          ),
      .I1      (in[129]              ),
      .I0      (out[129]             ),
      .O       (in[128]                )
   );
   (* BEL="X1/Y17/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut129 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[129]      ),
      .O       (out[130]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y17/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut129 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[130]          ),
      .I1      (in[130]              ),
      .I0      (out[130]             ),
      .O       (in[129]                )
   );
   (* BEL="X1/Y17/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut130 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[130]      ),
      .O       (out[131]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y17/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut130 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[131]          ),
      .I1      (in[131]              ),
      .I0      (out[131]             ),
      .O       (in[130]                )
   );
   (* BEL="X1/Y17/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut131 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[131]      ),
      .O       (out[132]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y17/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut131 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[132]          ),
      .I1      (in[132]              ),
      .I0      (out[132]             ),
      .O       (in[131]                )
   );
   (* BEL="X1/Y17/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut132 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[132]      ),
      .O       (out[133]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y17/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut132 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[133]          ),
      .I1      (in[133]              ),
      .I0      (out[133]             ),
      .O       (in[132]                )
   );
   (* BEL="X1/Y17/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut133 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[133]      ),
      .O       (out[134]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y17/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut133 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[134]          ),
      .I1      (in[134]              ),
      .I0      (out[134]             ),
      .O       (in[133]                )
   );
   (* BEL="X1/Y17/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut134 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[134]      ),
      .O       (out[135]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y17/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut134 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[135]          ),
      .I1      (in[135]              ),
      .I0      (out[135]             ),
      .O       (in[134]                )
   );
   (* BEL="X1/Y17/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut135 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[135]      ),
      .O       (out[136]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y17/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut135 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[136]          ),
      .I1      (in[136]              ),
      .I0      (out[136]             ),
      .O       (in[135]                )
   );
   (* BEL="X1/Y18/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut136 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[136]      ),
      .O       (out[137]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y18/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut136 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[137]          ),
      .I1      (in[137]              ),
      .I0      (out[137]             ),
      .O       (in[136]                )
   );
   (* BEL="X1/Y18/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut137 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[137]      ),
      .O       (out[138]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y18/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut137 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[138]          ),
      .I1      (in[138]              ),
      .I0      (out[138]             ),
      .O       (in[137]                )
   );
   (* BEL="X1/Y18/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut138 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[138]      ),
      .O       (out[139]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y18/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut138 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[139]          ),
      .I1      (in[139]              ),
      .I0      (out[139]             ),
      .O       (in[138]                )
   );
   (* BEL="X1/Y18/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut139 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[139]      ),
      .O       (out[140]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y18/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut139 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[140]          ),
      .I1      (in[140]              ),
      .I0      (out[140]             ),
      .O       (in[139]                )
   );
   (* BEL="X1/Y18/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut140 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[140]      ),
      .O       (out[141]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y18/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut140 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[141]          ),
      .I1      (in[141]              ),
      .I0      (out[141]             ),
      .O       (in[140]                )
   );
   (* BEL="X1/Y18/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut141 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[141]      ),
      .O       (out[142]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y18/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut141 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[142]          ),
      .I1      (in[142]              ),
      .I0      (out[142]             ),
      .O       (in[141]                )
   );
   (* BEL="X1/Y18/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut142 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[142]      ),
      .O       (out[143]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y18/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut142 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[143]          ),
      .I1      (in[143]              ),
      .I0      (out[143]             ),
      .O       (in[142]                )
   );
   (* BEL="X1/Y18/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut143 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[143]      ),
      .O       (out[144]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y18/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut143 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[144]          ),
      .I1      (in[144]              ),
      .I0      (out[144]             ),
      .O       (in[143]                )
   );
   (* BEL="X1/Y19/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut144 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[144]      ),
      .O       (out[145]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y19/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut144 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[145]          ),
      .I1      (in[145]              ),
      .I0      (out[145]             ),
      .O       (in[144]                )
   );
   (* BEL="X1/Y19/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut145 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[145]      ),
      .O       (out[146]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y19/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut145 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[146]          ),
      .I1      (in[146]              ),
      .I0      (out[146]             ),
      .O       (in[145]                )
   );
   (* BEL="X1/Y19/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut146 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[146]      ),
      .O       (out[147]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y19/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut146 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[147]          ),
      .I1      (in[147]              ),
      .I0      (out[147]             ),
      .O       (in[146]                )
   );
   (* BEL="X1/Y19/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut147 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[147]      ),
      .O       (out[148]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y19/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut147 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[148]          ),
      .I1      (in[148]              ),
      .I0      (out[148]             ),
      .O       (in[147]                )
   );
   (* BEL="X1/Y19/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut148 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[148]      ),
      .O       (out[149]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y19/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut148 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[149]          ),
      .I1      (in[149]              ),
      .I0      (out[149]             ),
      .O       (in[148]                )
   );
   (* BEL="X1/Y19/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut149 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[149]      ),
      .O       (out[150]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y19/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut149 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[150]          ),
      .I1      (in[150]              ),
      .I0      (out[150]             ),
      .O       (in[149]                )
   );
   (* BEL="X1/Y19/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut150 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[150]      ),
      .O       (out[151]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y19/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut150 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[151]          ),
      .I1      (in[151]              ),
      .I0      (out[151]             ),
      .O       (in[150]                )
   );
   (* BEL="X1/Y19/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut151 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[151]      ),
      .O       (out[152]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y19/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut151 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[152]          ),
      .I1      (in[152]              ),
      .I0      (out[152]             ),
      .O       (in[151]                )
   );
   (* BEL="X1/Y20/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut152 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[152]      ),
      .O       (out[153]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y20/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut152 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[153]          ),
      .I1      (in[153]              ),
      .I0      (out[153]             ),
      .O       (in[152]                )
   );
   (* BEL="X1/Y20/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut153 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[153]      ),
      .O       (out[154]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y20/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut153 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[154]          ),
      .I1      (in[154]              ),
      .I0      (out[154]             ),
      .O       (in[153]                )
   );
   (* BEL="X1/Y20/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut154 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[154]      ),
      .O       (out[155]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y20/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut154 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[155]          ),
      .I1      (in[155]              ),
      .I0      (out[155]             ),
      .O       (in[154]                )
   );
   (* BEL="X1/Y20/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut155 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[155]      ),
      .O       (out[156]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y20/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut155 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[156]          ),
      .I1      (in[156]              ),
      .I0      (out[156]             ),
      .O       (in[155]                )
   );
   (* BEL="X1/Y20/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut156 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[156]      ),
      .O       (out[157]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y20/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut156 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[157]          ),
      .I1      (in[157]              ),
      .I0      (out[157]             ),
      .O       (in[156]                )
   );
   (* BEL="X1/Y20/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut157 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[157]      ),
      .O       (out[158]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y20/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut157 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[158]          ),
      .I1      (in[158]              ),
      .I0      (out[158]             ),
      .O       (in[157]                )
   );
   (* BEL="X1/Y20/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut158 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[158]      ),
      .O       (out[159]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y20/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut158 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[159]          ),
      .I1      (in[159]              ),
      .I0      (out[159]             ),
      .O       (in[158]                )
   );
   (* BEL="X1/Y20/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut159 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[159]      ),
      .O       (out[160]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y20/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut159 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[160]          ),
      .I1      (in[160]              ),
      .I0      (out[160]             ),
      .O       (in[159]                )
   );
   (* BEL="X1/Y21/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut160 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[160]      ),
      .O       (out[161]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y21/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut160 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[161]          ),
      .I1      (in[161]              ),
      .I0      (out[161]             ),
      .O       (in[160]                )
   );
   (* BEL="X1/Y21/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut161 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[161]      ),
      .O       (out[162]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y21/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut161 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[162]          ),
      .I1      (in[162]              ),
      .I0      (out[162]             ),
      .O       (in[161]                )
   );
   (* BEL="X1/Y21/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut162 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[162]      ),
      .O       (out[163]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y21/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut162 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[163]          ),
      .I1      (in[163]              ),
      .I0      (out[163]             ),
      .O       (in[162]                )
   );
   (* BEL="X1/Y21/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut163 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[163]      ),
      .O       (out[164]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y21/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut163 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[164]          ),
      .I1      (in[164]              ),
      .I0      (out[164]             ),
      .O       (in[163]                )
   );
   (* BEL="X1/Y21/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut164 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[164]      ),
      .O       (out[165]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y21/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut164 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[165]          ),
      .I1      (in[165]              ),
      .I0      (out[165]             ),
      .O       (in[164]                )
   );
   (* BEL="X1/Y21/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut165 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[165]      ),
      .O       (out[166]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y21/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut165 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[166]          ),
      .I1      (in[166]              ),
      .I0      (out[166]             ),
      .O       (in[165]                )
   );
   (* BEL="X1/Y21/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut166 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[166]      ),
      .O       (out[167]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y21/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut166 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[167]          ),
      .I1      (in[167]              ),
      .I0      (out[167]             ),
      .O       (in[166]                )
   );
   (* BEL="X1/Y21/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut167 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[167]      ),
      .O       (out[168]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y21/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut167 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[168]          ),
      .I1      (in[168]              ),
      .I0      (out[168]             ),
      .O       (in[167]                )
   );
   (* BEL="X1/Y22/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut168 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[168]      ),
      .O       (out[169]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y22/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut168 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[169]          ),
      .I1      (in[169]              ),
      .I0      (out[169]             ),
      .O       (in[168]                )
   );
   (* BEL="X1/Y22/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut169 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[169]      ),
      .O       (out[170]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y22/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut169 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[170]          ),
      .I1      (in[170]              ),
      .I0      (out[170]             ),
      .O       (in[169]                )
   );
   (* BEL="X1/Y22/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut170 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[170]      ),
      .O       (out[171]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y22/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut170 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[171]          ),
      .I1      (in[171]              ),
      .I0      (out[171]             ),
      .O       (in[170]                )
   );
   (* BEL="X1/Y22/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut171 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[171]      ),
      .O       (out[172]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y22/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut171 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[172]          ),
      .I1      (in[172]              ),
      .I0      (out[172]             ),
      .O       (in[171]                )
   );
   (* BEL="X1/Y22/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut172 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[172]      ),
      .O       (out[173]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y22/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut172 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[173]          ),
      .I1      (in[173]              ),
      .I0      (out[173]             ),
      .O       (in[172]                )
   );
   (* BEL="X1/Y22/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut173 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[173]      ),
      .O       (out[174]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y22/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut173 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[174]          ),
      .I1      (in[174]              ),
      .I0      (out[174]             ),
      .O       (in[173]                )
   );
   (* BEL="X1/Y22/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut174 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[174]      ),
      .O       (out[175]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y22/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut174 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[175]          ),
      .I1      (in[175]              ),
      .I0      (out[175]             ),
      .O       (in[174]                )
   );
   (* BEL="X1/Y22/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut175 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[175]      ),
      .O       (out[176]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y22/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut175 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[176]          ),
      .I1      (in[176]              ),
      .I0      (out[176]             ),
      .O       (in[175]                )
   );
   (* BEL="X1/Y23/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut176 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[176]      ),
      .O       (out[177]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y23/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut176 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[177]          ),
      .I1      (in[177]              ),
      .I0      (out[177]             ),
      .O       (in[176]                )
   );
   (* BEL="X1/Y23/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut177 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[177]      ),
      .O       (out[178]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y23/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut177 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[178]          ),
      .I1      (in[178]              ),
      .I0      (out[178]             ),
      .O       (in[177]                )
   );
   (* BEL="X1/Y23/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut178 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[178]      ),
      .O       (out[179]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y23/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut178 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[179]          ),
      .I1      (in[179]              ),
      .I0      (out[179]             ),
      .O       (in[178]                )
   );
   (* BEL="X1/Y23/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut179 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[179]      ),
      .O       (out[180]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y23/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut179 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[180]          ),
      .I1      (in[180]              ),
      .I0      (out[180]             ),
      .O       (in[179]                )
   );
   (* BEL="X1/Y23/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut180 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[180]      ),
      .O       (out[181]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y23/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut180 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[181]          ),
      .I1      (in[181]              ),
      .I0      (out[181]             ),
      .O       (in[180]                )
   );
   (* BEL="X1/Y23/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut181 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[181]      ),
      .O       (out[182]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y23/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut181 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[182]          ),
      .I1      (in[182]              ),
      .I0      (out[182]             ),
      .O       (in[181]                )
   );
   (* BEL="X1/Y23/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut182 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[182]      ),
      .O       (out[183]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y23/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut182 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[183]          ),
      .I1      (in[183]              ),
      .I0      (out[183]             ),
      .O       (in[182]                )
   );
   (* BEL="X1/Y23/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut183 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[183]      ),
      .O       (out[184]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y23/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut183 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[184]          ),
      .I1      (in[184]              ),
      .I0      (out[184]             ),
      .O       (in[183]                )
   );
   (* BEL="X1/Y24/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut184 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[184]      ),
      .O       (out[185]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y24/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut184 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[185]          ),
      .I1      (in[185]              ),
      .I0      (out[185]             ),
      .O       (in[184]                )
   );
   (* BEL="X1/Y24/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut185 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[185]      ),
      .O       (out[186]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y24/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut185 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[186]          ),
      .I1      (in[186]              ),
      .I0      (out[186]             ),
      .O       (in[185]                )
   );
   (* BEL="X1/Y24/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut186 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[186]      ),
      .O       (out[187]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y24/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut186 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[187]          ),
      .I1      (in[187]              ),
      .I0      (out[187]             ),
      .O       (in[186]                )
   );
   (* BEL="X1/Y24/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut187 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[187]      ),
      .O       (out[188]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y24/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut187 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[188]          ),
      .I1      (in[188]              ),
      .I0      (out[188]             ),
      .O       (in[187]                )
   );
   (* BEL="X1/Y24/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut188 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[188]      ),
      .O       (out[189]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y24/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut188 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[189]          ),
      .I1      (in[189]              ),
      .I0      (out[189]             ),
      .O       (in[188]                )
   );
   (* BEL="X1/Y24/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut189 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[189]      ),
      .O       (out[190]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y24/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut189 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[190]          ),
      .I1      (in[190]              ),
      .I0      (out[190]             ),
      .O       (in[189]                )
   );
   (* BEL="X1/Y24/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut190 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[190]      ),
      .O       (out[191]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y24/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut190 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[191]          ),
      .I1      (in[191]              ),
      .I0      (out[191]             ),
      .O       (in[190]                )
   );
   (* BEL="X1/Y24/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut191 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[191]      ),
      .O       (out[192]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y24/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut191 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[192]          ),
      .I1      (in[192]              ),
      .I0      (out[192]             ),
      .O       (in[191]                )
   );
   (* BEL="X1/Y25/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut192 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[192]      ),
      .O       (out[193]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y25/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut192 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[193]          ),
      .I1      (in[193]              ),
      .I0      (out[193]             ),
      .O       (in[192]                )
   );
   (* BEL="X1/Y25/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut193 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[193]      ),
      .O       (out[194]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y25/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut193 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[194]          ),
      .I1      (in[194]              ),
      .I0      (out[194]             ),
      .O       (in[193]                )
   );
   (* BEL="X1/Y25/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut194 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[194]      ),
      .O       (out[195]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y25/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut194 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[195]          ),
      .I1      (in[195]              ),
      .I0      (out[195]             ),
      .O       (in[194]                )
   );
   (* BEL="X1/Y25/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut195 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[195]      ),
      .O       (out[196]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y25/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut195 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[196]          ),
      .I1      (in[196]              ),
      .I0      (out[196]             ),
      .O       (in[195]                )
   );
   (* BEL="X1/Y25/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut196 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[196]      ),
      .O       (out[197]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y25/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut196 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[197]          ),
      .I1      (in[197]              ),
      .I0      (out[197]             ),
      .O       (in[196]                )
   );
   (* BEL="X1/Y25/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut197 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[197]      ),
      .O       (out[198]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y25/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut197 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[198]          ),
      .I1      (in[198]              ),
      .I0      (out[198]             ),
      .O       (in[197]                )
   );
   (* BEL="X1/Y25/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut198 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[198]      ),
      .O       (out[199]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y25/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut198 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[199]          ),
      .I1      (in[199]              ),
      .I0      (out[199]             ),
      .O       (in[198]                )
   );
   (* BEL="X1/Y25/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut199 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[199]      ),
      .O       (out[200]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y25/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut199 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[200]          ),
      .I1      (in[200]              ),
      .I0      (out[200]             ),
      .O       (in[199]                )
   );
   (* BEL="X1/Y26/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut200 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[200]      ),
      .O       (out[201]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y26/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut200 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[201]          ),
      .I1      (in[201]              ),
      .I0      (out[201]             ),
      .O       (in[200]                )
   );
   (* BEL="X1/Y26/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut201 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[201]      ),
      .O       (out[202]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y26/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut201 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[202]          ),
      .I1      (in[202]              ),
      .I0      (out[202]             ),
      .O       (in[201]                )
   );
   (* BEL="X1/Y26/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut202 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[202]      ),
      .O       (out[203]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y26/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut202 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[203]          ),
      .I1      (in[203]              ),
      .I0      (out[203]             ),
      .O       (in[202]                )
   );
   (* BEL="X1/Y26/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut203 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[203]      ),
      .O       (out[204]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y26/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut203 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[204]          ),
      .I1      (in[204]              ),
      .I0      (out[204]             ),
      .O       (in[203]                )
   );
   (* BEL="X1/Y26/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut204 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[204]      ),
      .O       (out[205]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y26/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut204 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[205]          ),
      .I1      (in[205]              ),
      .I0      (out[205]             ),
      .O       (in[204]                )
   );
   (* BEL="X1/Y26/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut205 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[205]      ),
      .O       (out[206]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y26/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut205 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[206]          ),
      .I1      (in[206]              ),
      .I0      (out[206]             ),
      .O       (in[205]                )
   );
   (* BEL="X1/Y26/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut206 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[206]      ),
      .O       (out[207]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y26/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut206 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[207]          ),
      .I1      (in[207]              ),
      .I0      (out[207]             ),
      .O       (in[206]                )
   );
   (* BEL="X1/Y26/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut207 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[207]      ),
      .O       (out[208]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y26/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut207 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[208]          ),
      .I1      (in[208]              ),
      .I0      (out[208]             ),
      .O       (in[207]                )
   );
   (* BEL="X1/Y27/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut208 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[208]      ),
      .O       (out[209]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y27/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut208 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[209]          ),
      .I1      (in[209]              ),
      .I0      (out[209]             ),
      .O       (in[208]                )
   );
   (* BEL="X1/Y27/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut209 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[209]      ),
      .O       (out[210]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y27/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut209 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[210]          ),
      .I1      (in[210]              ),
      .I0      (out[210]             ),
      .O       (in[209]                )
   );
   (* BEL="X1/Y27/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut210 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[210]      ),
      .O       (out[211]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y27/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut210 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[211]          ),
      .I1      (in[211]              ),
      .I0      (out[211]             ),
      .O       (in[210]                )
   );
   (* BEL="X1/Y27/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut211 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[211]      ),
      .O       (out[212]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y27/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut211 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[212]          ),
      .I1      (in[212]              ),
      .I0      (out[212]             ),
      .O       (in[211]                )
   );
   (* BEL="X1/Y27/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut212 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[212]      ),
      .O       (out[213]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y27/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut212 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[213]          ),
      .I1      (in[213]              ),
      .I0      (out[213]             ),
      .O       (in[212]                )
   );
   (* BEL="X1/Y27/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut213 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[213]      ),
      .O       (out[214]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y27/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut213 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[214]          ),
      .I1      (in[214]              ),
      .I0      (out[214]             ),
      .O       (in[213]                )
   );
   (* BEL="X1/Y27/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut214 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[214]      ),
      .O       (out[215]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y27/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut214 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[215]          ),
      .I1      (in[215]              ),
      .I0      (out[215]             ),
      .O       (in[214]                )
   );
   (* BEL="X1/Y27/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut215 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[215]      ),
      .O       (out[216]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y27/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut215 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[216]          ),
      .I1      (in[216]              ),
      .I0      (out[216]             ),
      .O       (in[215]                )
   );
   (* BEL="X1/Y28/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut216 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[216]      ),
      .O       (out[217]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y28/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut216 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[217]          ),
      .I1      (in[217]              ),
      .I0      (out[217]             ),
      .O       (in[216]                )
   );
   (* BEL="X1/Y28/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut217 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[217]      ),
      .O       (out[218]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y28/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut217 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[218]          ),
      .I1      (in[218]              ),
      .I0      (out[218]             ),
      .O       (in[217]                )
   );
   (* BEL="X1/Y28/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut218 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[218]      ),
      .O       (out[219]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y28/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut218 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[219]          ),
      .I1      (in[219]              ),
      .I0      (out[219]             ),
      .O       (in[218]                )
   );
   (* BEL="X1/Y28/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut219 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[219]      ),
      .O       (out[220]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y28/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut219 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[220]          ),
      .I1      (in[220]              ),
      .I0      (out[220]             ),
      .O       (in[219]                )
   );
   (* BEL="X1/Y28/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut220 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[220]      ),
      .O       (out[221]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y28/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut220 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[221]          ),
      .I1      (in[221]              ),
      .I0      (out[221]             ),
      .O       (in[220]                )
   );
   (* BEL="X1/Y28/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut221 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[221]      ),
      .O       (out[222]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y28/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut221 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[222]          ),
      .I1      (in[222]              ),
      .I0      (out[222]             ),
      .O       (in[221]                )
   );
   (* BEL="X1/Y28/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut222 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[222]      ),
      .O       (out[223]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y28/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut222 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[223]          ),
      .I1      (in[223]              ),
      .I0      (out[223]             ),
      .O       (in[222]                )
   );
   (* BEL="X1/Y28/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut223 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[223]      ),
      .O       (out[224]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y28/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut223 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[224]          ),
      .I1      (in[224]              ),
      .I0      (out[224]             ),
      .O       (in[223]                )
   );
   (* BEL="X1/Y29/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut224 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[224]      ),
      .O       (out[225]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y29/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut224 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[225]          ),
      .I1      (in[225]              ),
      .I0      (out[225]             ),
      .O       (in[224]                )
   );
   (* BEL="X1/Y29/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut225 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[225]      ),
      .O       (out[226]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y29/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut225 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[226]          ),
      .I1      (in[226]              ),
      .I0      (out[226]             ),
      .O       (in[225]                )
   );
   (* BEL="X1/Y29/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut226 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[226]      ),
      .O       (out[227]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y29/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut226 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[227]          ),
      .I1      (in[227]              ),
      .I0      (out[227]             ),
      .O       (in[226]                )
   );
   (* BEL="X1/Y29/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut227 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[227]      ),
      .O       (out[228]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y29/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut227 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[228]          ),
      .I1      (in[228]              ),
      .I0      (out[228]             ),
      .O       (in[227]                )
   );
   (* BEL="X1/Y29/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut228 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[228]      ),
      .O       (out[229]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y29/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut228 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[229]          ),
      .I1      (in[229]              ),
      .I0      (out[229]             ),
      .O       (in[228]                )
   );
   (* BEL="X1/Y29/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut229 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[229]      ),
      .O       (out[230]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y29/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut229 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[230]          ),
      .I1      (in[230]              ),
      .I0      (out[230]             ),
      .O       (in[229]                )
   );
   (* BEL="X1/Y29/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut230 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[230]      ),
      .O       (out[231]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y29/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut230 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[231]          ),
      .I1      (in[231]              ),
      .I0      (out[231]             ),
      .O       (in[230]                )
   );
   (* BEL="X1/Y29/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut231 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[231]      ),
      .O       (out[232]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y29/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut231 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[232]          ),
      .I1      (in[232]              ),
      .I0      (out[232]             ),
      .O       (in[231]                )
   );
   (* BEL="X1/Y30/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut232 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[232]      ),
      .O       (out[233]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y30/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut232 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[233]          ),
      .I1      (in[233]              ),
      .I0      (out[233]             ),
      .O       (in[232]                )
   );
   (* BEL="X1/Y30/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut233 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[233]      ),
      .O       (out[234]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y30/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut233 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[234]          ),
      .I1      (in[234]              ),
      .I0      (out[234]             ),
      .O       (in[233]                )
   );
   (* BEL="X1/Y30/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut234 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[234]      ),
      .O       (out[235]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y30/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut234 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[235]          ),
      .I1      (in[235]              ),
      .I0      (out[235]             ),
      .O       (in[234]                )
   );
   (* BEL="X1/Y30/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut235 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[235]      ),
      .O       (out[236]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y30/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut235 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[236]          ),
      .I1      (in[236]              ),
      .I0      (out[236]             ),
      .O       (in[235]                )
   );
   (* BEL="X1/Y30/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut236 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[236]      ),
      .O       (out[237]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y30/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut236 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[237]          ),
      .I1      (in[237]              ),
      .I0      (out[237]             ),
      .O       (in[236]                )
   );
   (* BEL="X1/Y30/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut237 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[237]      ),
      .O       (out[238]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y30/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut237 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[238]          ),
      .I1      (in[238]              ),
      .I0      (out[238]             ),
      .O       (in[237]                )
   );
   (* BEL="X1/Y30/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut238 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[238]      ),
      .O       (out[239]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y30/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut238 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[239]          ),
      .I1      (in[239]              ),
      .I0      (out[239]             ),
      .O       (in[238]                )
   );
   (* BEL="X1/Y30/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut239 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[239]      ),
      .O       (out[240]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y30/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut239 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[240]          ),
      .I1      (in[240]              ),
      .I0      (out[240]             ),
      .O       (in[239]                )
   );
   (* BEL="X1/Y31/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut240 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[240]      ),
      .O       (out[241]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y31/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut240 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[241]          ),
      .I1      (in[241]              ),
      .I0      (out[241]             ),
      .O       (in[240]                )
   );
   (* BEL="X1/Y31/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut241 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[241]      ),
      .O       (out[242]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y31/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut241 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[242]          ),
      .I1      (in[242]              ),
      .I0      (out[242]             ),
      .O       (in[241]                )
   );
   (* BEL="X1/Y31/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut242 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[242]      ),
      .O       (out[243]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y31/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut242 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[243]          ),
      .I1      (in[243]              ),
      .I0      (out[243]             ),
      .O       (in[242]                )
   );
   (* BEL="X1/Y31/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut243 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[243]      ),
      .O       (out[244]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y31/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut243 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[244]          ),
      .I1      (in[244]              ),
      .I0      (out[244]             ),
      .O       (in[243]                )
   );
   (* BEL="X1/Y31/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut244 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[244]      ),
      .O       (out[245]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y31/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut244 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[245]          ),
      .I1      (in[245]              ),
      .I0      (out[245]             ),
      .O       (in[244]                )
   );
   (* BEL="X1/Y31/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut245 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[245]      ),
      .O       (out[246]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y31/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut245 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[246]          ),
      .I1      (in[246]              ),
      .I0      (out[246]             ),
      .O       (in[245]                )
   );
   (* BEL="X1/Y31/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut246 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[246]      ),
      .O       (out[247]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y31/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut246 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[247]          ),
      .I1      (in[247]              ),
      .I0      (out[247]             ),
      .O       (in[246]                )
   );
   (* BEL="X1/Y31/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut247 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[247]      ),
      .O       (out[248]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y31/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut247 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[248]          ),
      .I1      (in[248]              ),
      .I0      (out[248]             ),
      .O       (in[247]                )
   );
   (* BEL="X1/Y32/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut248 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[248]      ),
      .O       (out[249]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y32/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut248 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[249]          ),
      .I1      (in[249]              ),
      .I0      (out[249]             ),
      .O       (in[248]                )
   );
   (* BEL="X1/Y32/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut249 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[249]      ),
      .O       (out[250]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y32/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut249 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[250]          ),
      .I1      (in[250]              ),
      .I0      (out[250]             ),
      .O       (in[249]                )
   );
   (* BEL="X1/Y32/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut250 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[250]      ),
      .O       (out[251]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y32/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut250 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[251]          ),
      .I1      (in[251]              ),
      .I0      (out[251]             ),
      .O       (in[250]                )
   );
   (* BEL="X1/Y32/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut251 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[251]      ),
      .O       (out[252]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y32/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut251 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[252]          ),
      .I1      (in[252]              ),
      .I0      (out[252]             ),
      .O       (in[251]                )
   );
   (* BEL="X1/Y32/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut252 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[252]      ),
      .O       (out[253]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y32/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut252 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[253]          ),
      .I1      (in[253]              ),
      .I0      (out[253]             ),
      .O       (in[252]                )
   );
   (* BEL="X1/Y32/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut253 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[253]      ),
      .O       (out[254]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y32/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut253 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[254]          ),
      .I1      (in[254]              ),
      .I0      (out[254]             ),
      .O       (in[253]                )
   );
   (* BEL="X1/Y32/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut254 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[254]      ),
      .O       (out[255]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y32/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut254 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[255]          ),
      .I1      (in[255]              ),
      .I0      (out[255]             ),
      .O       (in[254]                )
   );
   (* BEL="X1/Y32/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) u_out_lut255 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (out[255]      ),
      .O       (out[256]    )
   );

   // i_ctrl   in[i+1]   out[i+1]  |  in[i]
   // ---------------------------------------
   //    0       0          0      |   0 
   //    0       0          1      |   0 
   //    0       1          0      |   1 
   //    0       1          1      |   1 
   //    1       0          0      |   0 
   //    1       0          1      |   1 
   //    1       1          0      |   0 
   //    1       1          1      |   1 

   (* BEL="X2/Y32/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'b0000000010101100   )
   ) u_in_lut255 (
      .I3      (1'b0                   ),
      .I2      (i_ctrl[256]          ),
      .I1      (in[256]              ),
      .I0      (out[256]             ),
      .O       (in[255]                )
   );

assign o_dl = in[0];

endmodule

