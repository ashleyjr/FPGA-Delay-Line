module x_delay_line (
   input    logic                         i_clk,
   input    logic                         i_dl,
   output   logic [256-1:0]          o_data
);

logic [256:0]   p0_dl;
logic [256-1:0] p1_dl;
logic [256-1:0] p2_dl;

assign p0_dl[0] = i_dl;

   (* BEL="X9/Y1/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut0 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[0]    ),
      .O       (p0_dl[1]  )
   );

   (* BEL="X9/Y1/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut1 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[1]    ),
      .O       (p0_dl[2]  )
   );

   (* BEL="X9/Y1/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut2 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[2]    ),
      .O       (p0_dl[3]  )
   );

   (* BEL="X9/Y1/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut3 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[3]    ),
      .O       (p0_dl[4]  )
   );

   (* BEL="X9/Y1/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut4 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[4]    ),
      .O       (p0_dl[5]  )
   );

   (* BEL="X9/Y1/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut5 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[5]    ),
      .O       (p0_dl[6]  )
   );

   (* BEL="X9/Y1/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut6 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[6]    ),
      .O       (p0_dl[7]  )
   );

   (* BEL="X9/Y1/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut7 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[7]    ),
      .O       (p0_dl[8]  )
   );

   (* BEL="X9/Y2/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut8 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[8]    ),
      .O       (p0_dl[9]  )
   );

   (* BEL="X9/Y2/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut9 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[9]    ),
      .O       (p0_dl[10]  )
   );

   (* BEL="X9/Y2/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut10 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[10]    ),
      .O       (p0_dl[11]  )
   );

   (* BEL="X9/Y2/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut11 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[11]    ),
      .O       (p0_dl[12]  )
   );

   (* BEL="X9/Y2/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut12 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[12]    ),
      .O       (p0_dl[13]  )
   );

   (* BEL="X9/Y2/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut13 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[13]    ),
      .O       (p0_dl[14]  )
   );

   (* BEL="X9/Y2/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut14 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[14]    ),
      .O       (p0_dl[15]  )
   );

   (* BEL="X9/Y2/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut15 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[15]    ),
      .O       (p0_dl[16]  )
   );

   (* BEL="X9/Y3/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut16 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[16]    ),
      .O       (p0_dl[17]  )
   );

   (* BEL="X9/Y3/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut17 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[17]    ),
      .O       (p0_dl[18]  )
   );

   (* BEL="X9/Y3/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut18 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[18]    ),
      .O       (p0_dl[19]  )
   );

   (* BEL="X9/Y3/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut19 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[19]    ),
      .O       (p0_dl[20]  )
   );

   (* BEL="X9/Y3/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut20 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[20]    ),
      .O       (p0_dl[21]  )
   );

   (* BEL="X9/Y3/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut21 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[21]    ),
      .O       (p0_dl[22]  )
   );

   (* BEL="X9/Y3/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut22 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[22]    ),
      .O       (p0_dl[23]  )
   );

   (* BEL="X9/Y3/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut23 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[23]    ),
      .O       (p0_dl[24]  )
   );

   (* BEL="X9/Y4/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut24 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[24]    ),
      .O       (p0_dl[25]  )
   );

   (* BEL="X9/Y4/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut25 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[25]    ),
      .O       (p0_dl[26]  )
   );

   (* BEL="X9/Y4/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut26 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[26]    ),
      .O       (p0_dl[27]  )
   );

   (* BEL="X9/Y4/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut27 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[27]    ),
      .O       (p0_dl[28]  )
   );

   (* BEL="X9/Y4/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut28 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[28]    ),
      .O       (p0_dl[29]  )
   );

   (* BEL="X9/Y4/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut29 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[29]    ),
      .O       (p0_dl[30]  )
   );

   (* BEL="X9/Y4/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut30 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[30]    ),
      .O       (p0_dl[31]  )
   );

   (* BEL="X9/Y4/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut31 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[31]    ),
      .O       (p0_dl[32]  )
   );

   (* BEL="X9/Y5/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut32 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[32]    ),
      .O       (p0_dl[33]  )
   );

   (* BEL="X9/Y5/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut33 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[33]    ),
      .O       (p0_dl[34]  )
   );

   (* BEL="X9/Y5/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut34 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[34]    ),
      .O       (p0_dl[35]  )
   );

   (* BEL="X9/Y5/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut35 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[35]    ),
      .O       (p0_dl[36]  )
   );

   (* BEL="X9/Y5/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut36 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[36]    ),
      .O       (p0_dl[37]  )
   );

   (* BEL="X9/Y5/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut37 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[37]    ),
      .O       (p0_dl[38]  )
   );

   (* BEL="X9/Y5/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut38 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[38]    ),
      .O       (p0_dl[39]  )
   );

   (* BEL="X9/Y5/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut39 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[39]    ),
      .O       (p0_dl[40]  )
   );

   (* BEL="X9/Y6/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut40 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[40]    ),
      .O       (p0_dl[41]  )
   );

   (* BEL="X9/Y6/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut41 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[41]    ),
      .O       (p0_dl[42]  )
   );

   (* BEL="X9/Y6/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut42 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[42]    ),
      .O       (p0_dl[43]  )
   );

   (* BEL="X9/Y6/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut43 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[43]    ),
      .O       (p0_dl[44]  )
   );

   (* BEL="X9/Y6/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut44 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[44]    ),
      .O       (p0_dl[45]  )
   );

   (* BEL="X9/Y6/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut45 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[45]    ),
      .O       (p0_dl[46]  )
   );

   (* BEL="X9/Y6/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut46 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[46]    ),
      .O       (p0_dl[47]  )
   );

   (* BEL="X9/Y6/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut47 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[47]    ),
      .O       (p0_dl[48]  )
   );

   (* BEL="X9/Y7/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut48 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[48]    ),
      .O       (p0_dl[49]  )
   );

   (* BEL="X9/Y7/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut49 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[49]    ),
      .O       (p0_dl[50]  )
   );

   (* BEL="X9/Y7/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut50 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[50]    ),
      .O       (p0_dl[51]  )
   );

   (* BEL="X9/Y7/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut51 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[51]    ),
      .O       (p0_dl[52]  )
   );

   (* BEL="X9/Y7/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut52 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[52]    ),
      .O       (p0_dl[53]  )
   );

   (* BEL="X9/Y7/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut53 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[53]    ),
      .O       (p0_dl[54]  )
   );

   (* BEL="X9/Y7/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut54 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[54]    ),
      .O       (p0_dl[55]  )
   );

   (* BEL="X9/Y7/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut55 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[55]    ),
      .O       (p0_dl[56]  )
   );

   (* BEL="X9/Y8/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut56 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[56]    ),
      .O       (p0_dl[57]  )
   );

   (* BEL="X9/Y8/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut57 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[57]    ),
      .O       (p0_dl[58]  )
   );

   (* BEL="X9/Y8/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut58 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[58]    ),
      .O       (p0_dl[59]  )
   );

   (* BEL="X9/Y8/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut59 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[59]    ),
      .O       (p0_dl[60]  )
   );

   (* BEL="X9/Y8/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut60 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[60]    ),
      .O       (p0_dl[61]  )
   );

   (* BEL="X9/Y8/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut61 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[61]    ),
      .O       (p0_dl[62]  )
   );

   (* BEL="X9/Y8/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut62 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[62]    ),
      .O       (p0_dl[63]  )
   );

   (* BEL="X9/Y8/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut63 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[63]    ),
      .O       (p0_dl[64]  )
   );

   (* BEL="X9/Y9/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut64 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[64]    ),
      .O       (p0_dl[65]  )
   );

   (* BEL="X9/Y9/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut65 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[65]    ),
      .O       (p0_dl[66]  )
   );

   (* BEL="X9/Y9/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut66 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[66]    ),
      .O       (p0_dl[67]  )
   );

   (* BEL="X9/Y9/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut67 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[67]    ),
      .O       (p0_dl[68]  )
   );

   (* BEL="X9/Y9/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut68 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[68]    ),
      .O       (p0_dl[69]  )
   );

   (* BEL="X9/Y9/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut69 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[69]    ),
      .O       (p0_dl[70]  )
   );

   (* BEL="X9/Y9/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut70 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[70]    ),
      .O       (p0_dl[71]  )
   );

   (* BEL="X9/Y9/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut71 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[71]    ),
      .O       (p0_dl[72]  )
   );

   (* BEL="X9/Y10/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut72 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[72]    ),
      .O       (p0_dl[73]  )
   );

   (* BEL="X9/Y10/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut73 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[73]    ),
      .O       (p0_dl[74]  )
   );

   (* BEL="X9/Y10/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut74 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[74]    ),
      .O       (p0_dl[75]  )
   );

   (* BEL="X9/Y10/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut75 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[75]    ),
      .O       (p0_dl[76]  )
   );

   (* BEL="X9/Y10/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut76 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[76]    ),
      .O       (p0_dl[77]  )
   );

   (* BEL="X9/Y10/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut77 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[77]    ),
      .O       (p0_dl[78]  )
   );

   (* BEL="X9/Y10/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut78 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[78]    ),
      .O       (p0_dl[79]  )
   );

   (* BEL="X9/Y10/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut79 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[79]    ),
      .O       (p0_dl[80]  )
   );

   (* BEL="X9/Y11/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut80 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[80]    ),
      .O       (p0_dl[81]  )
   );

   (* BEL="X9/Y11/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut81 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[81]    ),
      .O       (p0_dl[82]  )
   );

   (* BEL="X9/Y11/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut82 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[82]    ),
      .O       (p0_dl[83]  )
   );

   (* BEL="X9/Y11/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut83 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[83]    ),
      .O       (p0_dl[84]  )
   );

   (* BEL="X9/Y11/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut84 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[84]    ),
      .O       (p0_dl[85]  )
   );

   (* BEL="X9/Y11/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut85 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[85]    ),
      .O       (p0_dl[86]  )
   );

   (* BEL="X9/Y11/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut86 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[86]    ),
      .O       (p0_dl[87]  )
   );

   (* BEL="X9/Y11/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut87 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[87]    ),
      .O       (p0_dl[88]  )
   );

   (* BEL="X9/Y12/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut88 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[88]    ),
      .O       (p0_dl[89]  )
   );

   (* BEL="X9/Y12/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut89 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[89]    ),
      .O       (p0_dl[90]  )
   );

   (* BEL="X9/Y12/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut90 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[90]    ),
      .O       (p0_dl[91]  )
   );

   (* BEL="X9/Y12/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut91 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[91]    ),
      .O       (p0_dl[92]  )
   );

   (* BEL="X9/Y12/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut92 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[92]    ),
      .O       (p0_dl[93]  )
   );

   (* BEL="X9/Y12/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut93 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[93]    ),
      .O       (p0_dl[94]  )
   );

   (* BEL="X9/Y12/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut94 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[94]    ),
      .O       (p0_dl[95]  )
   );

   (* BEL="X9/Y12/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut95 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[95]    ),
      .O       (p0_dl[96]  )
   );

   (* BEL="X9/Y13/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut96 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[96]    ),
      .O       (p0_dl[97]  )
   );

   (* BEL="X9/Y13/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut97 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[97]    ),
      .O       (p0_dl[98]  )
   );

   (* BEL="X9/Y13/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut98 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[98]    ),
      .O       (p0_dl[99]  )
   );

   (* BEL="X9/Y13/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut99 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[99]    ),
      .O       (p0_dl[100]  )
   );

   (* BEL="X9/Y13/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut100 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[100]    ),
      .O       (p0_dl[101]  )
   );

   (* BEL="X9/Y13/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut101 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[101]    ),
      .O       (p0_dl[102]  )
   );

   (* BEL="X9/Y13/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut102 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[102]    ),
      .O       (p0_dl[103]  )
   );

   (* BEL="X9/Y13/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut103 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[103]    ),
      .O       (p0_dl[104]  )
   );

   (* BEL="X9/Y14/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut104 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[104]    ),
      .O       (p0_dl[105]  )
   );

   (* BEL="X9/Y14/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut105 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[105]    ),
      .O       (p0_dl[106]  )
   );

   (* BEL="X9/Y14/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut106 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[106]    ),
      .O       (p0_dl[107]  )
   );

   (* BEL="X9/Y14/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut107 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[107]    ),
      .O       (p0_dl[108]  )
   );

   (* BEL="X9/Y14/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut108 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[108]    ),
      .O       (p0_dl[109]  )
   );

   (* BEL="X9/Y14/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut109 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[109]    ),
      .O       (p0_dl[110]  )
   );

   (* BEL="X9/Y14/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut110 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[110]    ),
      .O       (p0_dl[111]  )
   );

   (* BEL="X9/Y14/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut111 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[111]    ),
      .O       (p0_dl[112]  )
   );

   (* BEL="X9/Y15/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut112 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[112]    ),
      .O       (p0_dl[113]  )
   );

   (* BEL="X9/Y15/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut113 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[113]    ),
      .O       (p0_dl[114]  )
   );

   (* BEL="X9/Y15/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut114 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[114]    ),
      .O       (p0_dl[115]  )
   );

   (* BEL="X9/Y15/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut115 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[115]    ),
      .O       (p0_dl[116]  )
   );

   (* BEL="X9/Y15/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut116 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[116]    ),
      .O       (p0_dl[117]  )
   );

   (* BEL="X9/Y15/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut117 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[117]    ),
      .O       (p0_dl[118]  )
   );

   (* BEL="X9/Y15/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut118 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[118]    ),
      .O       (p0_dl[119]  )
   );

   (* BEL="X9/Y15/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut119 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[119]    ),
      .O       (p0_dl[120]  )
   );

   (* BEL="X9/Y16/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut120 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[120]    ),
      .O       (p0_dl[121]  )
   );

   (* BEL="X9/Y16/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut121 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[121]    ),
      .O       (p0_dl[122]  )
   );

   (* BEL="X9/Y16/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut122 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[122]    ),
      .O       (p0_dl[123]  )
   );

   (* BEL="X9/Y16/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut123 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[123]    ),
      .O       (p0_dl[124]  )
   );

   (* BEL="X9/Y16/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut124 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[124]    ),
      .O       (p0_dl[125]  )
   );

   (* BEL="X9/Y16/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut125 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[125]    ),
      .O       (p0_dl[126]  )
   );

   (* BEL="X9/Y16/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut126 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[126]    ),
      .O       (p0_dl[127]  )
   );

   (* BEL="X9/Y16/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut127 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[127]    ),
      .O       (p0_dl[128]  )
   );

   (* BEL="X9/Y17/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut128 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[128]    ),
      .O       (p0_dl[129]  )
   );

   (* BEL="X9/Y17/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut129 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[129]    ),
      .O       (p0_dl[130]  )
   );

   (* BEL="X9/Y17/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut130 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[130]    ),
      .O       (p0_dl[131]  )
   );

   (* BEL="X9/Y17/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut131 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[131]    ),
      .O       (p0_dl[132]  )
   );

   (* BEL="X9/Y17/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut132 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[132]    ),
      .O       (p0_dl[133]  )
   );

   (* BEL="X9/Y17/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut133 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[133]    ),
      .O       (p0_dl[134]  )
   );

   (* BEL="X9/Y17/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut134 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[134]    ),
      .O       (p0_dl[135]  )
   );

   (* BEL="X9/Y17/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut135 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[135]    ),
      .O       (p0_dl[136]  )
   );

   (* BEL="X9/Y18/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut136 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[136]    ),
      .O       (p0_dl[137]  )
   );

   (* BEL="X9/Y18/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut137 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[137]    ),
      .O       (p0_dl[138]  )
   );

   (* BEL="X9/Y18/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut138 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[138]    ),
      .O       (p0_dl[139]  )
   );

   (* BEL="X9/Y18/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut139 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[139]    ),
      .O       (p0_dl[140]  )
   );

   (* BEL="X9/Y18/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut140 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[140]    ),
      .O       (p0_dl[141]  )
   );

   (* BEL="X9/Y18/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut141 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[141]    ),
      .O       (p0_dl[142]  )
   );

   (* BEL="X9/Y18/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut142 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[142]    ),
      .O       (p0_dl[143]  )
   );

   (* BEL="X9/Y18/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut143 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[143]    ),
      .O       (p0_dl[144]  )
   );

   (* BEL="X9/Y19/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut144 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[144]    ),
      .O       (p0_dl[145]  )
   );

   (* BEL="X9/Y19/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut145 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[145]    ),
      .O       (p0_dl[146]  )
   );

   (* BEL="X9/Y19/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut146 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[146]    ),
      .O       (p0_dl[147]  )
   );

   (* BEL="X9/Y19/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut147 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[147]    ),
      .O       (p0_dl[148]  )
   );

   (* BEL="X9/Y19/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut148 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[148]    ),
      .O       (p0_dl[149]  )
   );

   (* BEL="X9/Y19/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut149 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[149]    ),
      .O       (p0_dl[150]  )
   );

   (* BEL="X9/Y19/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut150 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[150]    ),
      .O       (p0_dl[151]  )
   );

   (* BEL="X9/Y19/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut151 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[151]    ),
      .O       (p0_dl[152]  )
   );

   (* BEL="X9/Y20/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut152 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[152]    ),
      .O       (p0_dl[153]  )
   );

   (* BEL="X9/Y20/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut153 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[153]    ),
      .O       (p0_dl[154]  )
   );

   (* BEL="X9/Y20/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut154 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[154]    ),
      .O       (p0_dl[155]  )
   );

   (* BEL="X9/Y20/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut155 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[155]    ),
      .O       (p0_dl[156]  )
   );

   (* BEL="X9/Y20/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut156 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[156]    ),
      .O       (p0_dl[157]  )
   );

   (* BEL="X9/Y20/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut157 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[157]    ),
      .O       (p0_dl[158]  )
   );

   (* BEL="X9/Y20/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut158 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[158]    ),
      .O       (p0_dl[159]  )
   );

   (* BEL="X9/Y20/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut159 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[159]    ),
      .O       (p0_dl[160]  )
   );

   (* BEL="X9/Y21/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut160 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[160]    ),
      .O       (p0_dl[161]  )
   );

   (* BEL="X9/Y21/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut161 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[161]    ),
      .O       (p0_dl[162]  )
   );

   (* BEL="X9/Y21/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut162 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[162]    ),
      .O       (p0_dl[163]  )
   );

   (* BEL="X9/Y21/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut163 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[163]    ),
      .O       (p0_dl[164]  )
   );

   (* BEL="X9/Y21/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut164 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[164]    ),
      .O       (p0_dl[165]  )
   );

   (* BEL="X9/Y21/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut165 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[165]    ),
      .O       (p0_dl[166]  )
   );

   (* BEL="X9/Y21/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut166 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[166]    ),
      .O       (p0_dl[167]  )
   );

   (* BEL="X9/Y21/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut167 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[167]    ),
      .O       (p0_dl[168]  )
   );

   (* BEL="X9/Y22/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut168 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[168]    ),
      .O       (p0_dl[169]  )
   );

   (* BEL="X9/Y22/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut169 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[169]    ),
      .O       (p0_dl[170]  )
   );

   (* BEL="X9/Y22/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut170 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[170]    ),
      .O       (p0_dl[171]  )
   );

   (* BEL="X9/Y22/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut171 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[171]    ),
      .O       (p0_dl[172]  )
   );

   (* BEL="X9/Y22/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut172 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[172]    ),
      .O       (p0_dl[173]  )
   );

   (* BEL="X9/Y22/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut173 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[173]    ),
      .O       (p0_dl[174]  )
   );

   (* BEL="X9/Y22/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut174 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[174]    ),
      .O       (p0_dl[175]  )
   );

   (* BEL="X9/Y22/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut175 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[175]    ),
      .O       (p0_dl[176]  )
   );

   (* BEL="X9/Y23/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut176 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[176]    ),
      .O       (p0_dl[177]  )
   );

   (* BEL="X9/Y23/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut177 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[177]    ),
      .O       (p0_dl[178]  )
   );

   (* BEL="X9/Y23/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut178 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[178]    ),
      .O       (p0_dl[179]  )
   );

   (* BEL="X9/Y23/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut179 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[179]    ),
      .O       (p0_dl[180]  )
   );

   (* BEL="X9/Y23/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut180 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[180]    ),
      .O       (p0_dl[181]  )
   );

   (* BEL="X9/Y23/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut181 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[181]    ),
      .O       (p0_dl[182]  )
   );

   (* BEL="X9/Y23/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut182 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[182]    ),
      .O       (p0_dl[183]  )
   );

   (* BEL="X9/Y23/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut183 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[183]    ),
      .O       (p0_dl[184]  )
   );

   (* BEL="X9/Y24/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut184 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[184]    ),
      .O       (p0_dl[185]  )
   );

   (* BEL="X9/Y24/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut185 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[185]    ),
      .O       (p0_dl[186]  )
   );

   (* BEL="X9/Y24/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut186 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[186]    ),
      .O       (p0_dl[187]  )
   );

   (* BEL="X9/Y24/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut187 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[187]    ),
      .O       (p0_dl[188]  )
   );

   (* BEL="X9/Y24/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut188 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[188]    ),
      .O       (p0_dl[189]  )
   );

   (* BEL="X9/Y24/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut189 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[189]    ),
      .O       (p0_dl[190]  )
   );

   (* BEL="X9/Y24/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut190 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[190]    ),
      .O       (p0_dl[191]  )
   );

   (* BEL="X9/Y24/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut191 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[191]    ),
      .O       (p0_dl[192]  )
   );

   (* BEL="X9/Y25/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut192 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[192]    ),
      .O       (p0_dl[193]  )
   );

   (* BEL="X9/Y25/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut193 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[193]    ),
      .O       (p0_dl[194]  )
   );

   (* BEL="X9/Y25/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut194 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[194]    ),
      .O       (p0_dl[195]  )
   );

   (* BEL="X9/Y25/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut195 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[195]    ),
      .O       (p0_dl[196]  )
   );

   (* BEL="X9/Y25/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut196 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[196]    ),
      .O       (p0_dl[197]  )
   );

   (* BEL="X9/Y25/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut197 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[197]    ),
      .O       (p0_dl[198]  )
   );

   (* BEL="X9/Y25/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut198 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[198]    ),
      .O       (p0_dl[199]  )
   );

   (* BEL="X9/Y25/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut199 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[199]    ),
      .O       (p0_dl[200]  )
   );

   (* BEL="X9/Y26/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut200 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[200]    ),
      .O       (p0_dl[201]  )
   );

   (* BEL="X9/Y26/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut201 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[201]    ),
      .O       (p0_dl[202]  )
   );

   (* BEL="X9/Y26/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut202 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[202]    ),
      .O       (p0_dl[203]  )
   );

   (* BEL="X9/Y26/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut203 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[203]    ),
      .O       (p0_dl[204]  )
   );

   (* BEL="X9/Y26/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut204 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[204]    ),
      .O       (p0_dl[205]  )
   );

   (* BEL="X9/Y26/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut205 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[205]    ),
      .O       (p0_dl[206]  )
   );

   (* BEL="X9/Y26/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut206 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[206]    ),
      .O       (p0_dl[207]  )
   );

   (* BEL="X9/Y26/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut207 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[207]    ),
      .O       (p0_dl[208]  )
   );

   (* BEL="X9/Y27/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut208 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[208]    ),
      .O       (p0_dl[209]  )
   );

   (* BEL="X9/Y27/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut209 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[209]    ),
      .O       (p0_dl[210]  )
   );

   (* BEL="X9/Y27/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut210 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[210]    ),
      .O       (p0_dl[211]  )
   );

   (* BEL="X9/Y27/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut211 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[211]    ),
      .O       (p0_dl[212]  )
   );

   (* BEL="X9/Y27/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut212 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[212]    ),
      .O       (p0_dl[213]  )
   );

   (* BEL="X9/Y27/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut213 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[213]    ),
      .O       (p0_dl[214]  )
   );

   (* BEL="X9/Y27/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut214 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[214]    ),
      .O       (p0_dl[215]  )
   );

   (* BEL="X9/Y27/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut215 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[215]    ),
      .O       (p0_dl[216]  )
   );

   (* BEL="X9/Y28/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut216 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[216]    ),
      .O       (p0_dl[217]  )
   );

   (* BEL="X9/Y28/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut217 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[217]    ),
      .O       (p0_dl[218]  )
   );

   (* BEL="X9/Y28/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut218 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[218]    ),
      .O       (p0_dl[219]  )
   );

   (* BEL="X9/Y28/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut219 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[219]    ),
      .O       (p0_dl[220]  )
   );

   (* BEL="X9/Y28/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut220 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[220]    ),
      .O       (p0_dl[221]  )
   );

   (* BEL="X9/Y28/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut221 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[221]    ),
      .O       (p0_dl[222]  )
   );

   (* BEL="X9/Y28/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut222 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[222]    ),
      .O       (p0_dl[223]  )
   );

   (* BEL="X9/Y28/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut223 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[223]    ),
      .O       (p0_dl[224]  )
   );

   (* BEL="X9/Y29/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut224 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[224]    ),
      .O       (p0_dl[225]  )
   );

   (* BEL="X9/Y29/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut225 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[225]    ),
      .O       (p0_dl[226]  )
   );

   (* BEL="X9/Y29/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut226 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[226]    ),
      .O       (p0_dl[227]  )
   );

   (* BEL="X9/Y29/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut227 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[227]    ),
      .O       (p0_dl[228]  )
   );

   (* BEL="X9/Y29/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut228 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[228]    ),
      .O       (p0_dl[229]  )
   );

   (* BEL="X9/Y29/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut229 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[229]    ),
      .O       (p0_dl[230]  )
   );

   (* BEL="X9/Y29/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut230 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[230]    ),
      .O       (p0_dl[231]  )
   );

   (* BEL="X9/Y29/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut231 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[231]    ),
      .O       (p0_dl[232]  )
   );

   (* BEL="X9/Y30/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut232 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[232]    ),
      .O       (p0_dl[233]  )
   );

   (* BEL="X9/Y30/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut233 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[233]    ),
      .O       (p0_dl[234]  )
   );

   (* BEL="X9/Y30/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut234 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[234]    ),
      .O       (p0_dl[235]  )
   );

   (* BEL="X9/Y30/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut235 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[235]    ),
      .O       (p0_dl[236]  )
   );

   (* BEL="X9/Y30/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut236 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[236]    ),
      .O       (p0_dl[237]  )
   );

   (* BEL="X9/Y30/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut237 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[237]    ),
      .O       (p0_dl[238]  )
   );

   (* BEL="X9/Y30/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut238 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[238]    ),
      .O       (p0_dl[239]  )
   );

   (* BEL="X9/Y30/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut239 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[239]    ),
      .O       (p0_dl[240]  )
   );

   (* BEL="X9/Y31/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut240 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[240]    ),
      .O       (p0_dl[241]  )
   );

   (* BEL="X9/Y31/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut241 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[241]    ),
      .O       (p0_dl[242]  )
   );

   (* BEL="X9/Y31/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut242 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[242]    ),
      .O       (p0_dl[243]  )
   );

   (* BEL="X9/Y31/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut243 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[243]    ),
      .O       (p0_dl[244]  )
   );

   (* BEL="X9/Y31/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut244 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[244]    ),
      .O       (p0_dl[245]  )
   );

   (* BEL="X9/Y31/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut245 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[245]    ),
      .O       (p0_dl[246]  )
   );

   (* BEL="X9/Y31/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut246 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[246]    ),
      .O       (p0_dl[247]  )
   );

   (* BEL="X9/Y31/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut247 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[247]    ),
      .O       (p0_dl[248]  )
   );

   (* BEL="X9/Y32/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut248 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[248]    ),
      .O       (p0_dl[249]  )
   );

   (* BEL="X9/Y32/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut249 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[249]    ),
      .O       (p0_dl[250]  )
   );

   (* BEL="X9/Y32/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut250 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[250]    ),
      .O       (p0_dl[251]  )
   );

   (* BEL="X9/Y32/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut251 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[251]    ),
      .O       (p0_dl[252]  )
   );

   (* BEL="X9/Y32/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut252 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[252]    ),
      .O       (p0_dl[253]  )
   );

   (* BEL="X9/Y32/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut253 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[253]    ),
      .O       (p0_dl[254]  )
   );

   (* BEL="X9/Y32/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut254 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[254]    ),
      .O       (p0_dl[255]  )
   );

   (* BEL="X9/Y32/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut255 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[255]    ),
      .O       (p0_dl[256]  )
   );


   (* BEL="X10/Y1/lc0" *)
   SB_DFF  dff_2_0 (
      .C       (i_clk         ),
      .D       (p0_dl[1]  ),
      .Q       (p1_dl[0]    )
   );

   (* BEL="X11/Y1/lc0" *)
   SB_DFF  dff_3_0 (
      .C       (i_clk         ),
      .D       (p1_dl[0]    ),
      .Q       (o_data[0]   )
   );

   (* BEL="X10/Y1/lc1" *)
   SB_DFF  dff_2_1 (
      .C       (i_clk         ),
      .D       (p0_dl[2]  ),
      .Q       (p1_dl[1]    )
   );

   (* BEL="X11/Y1/lc1" *)
   SB_DFF  dff_3_1 (
      .C       (i_clk         ),
      .D       (p1_dl[1]    ),
      .Q       (o_data[1]   )
   );

   (* BEL="X10/Y1/lc2" *)
   SB_DFF  dff_2_2 (
      .C       (i_clk         ),
      .D       (p0_dl[3]  ),
      .Q       (p1_dl[2]    )
   );

   (* BEL="X11/Y1/lc2" *)
   SB_DFF  dff_3_2 (
      .C       (i_clk         ),
      .D       (p1_dl[2]    ),
      .Q       (o_data[2]   )
   );

   (* BEL="X10/Y1/lc3" *)
   SB_DFF  dff_2_3 (
      .C       (i_clk         ),
      .D       (p0_dl[4]  ),
      .Q       (p1_dl[3]    )
   );

   (* BEL="X11/Y1/lc3" *)
   SB_DFF  dff_3_3 (
      .C       (i_clk         ),
      .D       (p1_dl[3]    ),
      .Q       (o_data[3]   )
   );

   (* BEL="X10/Y1/lc4" *)
   SB_DFF  dff_2_4 (
      .C       (i_clk         ),
      .D       (p0_dl[5]  ),
      .Q       (p1_dl[4]    )
   );

   (* BEL="X11/Y1/lc4" *)
   SB_DFF  dff_3_4 (
      .C       (i_clk         ),
      .D       (p1_dl[4]    ),
      .Q       (o_data[4]   )
   );

   (* BEL="X10/Y1/lc5" *)
   SB_DFF  dff_2_5 (
      .C       (i_clk         ),
      .D       (p0_dl[6]  ),
      .Q       (p1_dl[5]    )
   );

   (* BEL="X11/Y1/lc5" *)
   SB_DFF  dff_3_5 (
      .C       (i_clk         ),
      .D       (p1_dl[5]    ),
      .Q       (o_data[5]   )
   );

   (* BEL="X10/Y1/lc6" *)
   SB_DFF  dff_2_6 (
      .C       (i_clk         ),
      .D       (p0_dl[7]  ),
      .Q       (p1_dl[6]    )
   );

   (* BEL="X11/Y1/lc6" *)
   SB_DFF  dff_3_6 (
      .C       (i_clk         ),
      .D       (p1_dl[6]    ),
      .Q       (o_data[6]   )
   );

   (* BEL="X10/Y1/lc7" *)
   SB_DFF  dff_2_7 (
      .C       (i_clk         ),
      .D       (p0_dl[8]  ),
      .Q       (p1_dl[7]    )
   );

   (* BEL="X11/Y1/lc7" *)
   SB_DFF  dff_3_7 (
      .C       (i_clk         ),
      .D       (p1_dl[7]    ),
      .Q       (o_data[7]   )
   );

   (* BEL="X10/Y2/lc0" *)
   SB_DFF  dff_2_8 (
      .C       (i_clk         ),
      .D       (p0_dl[9]  ),
      .Q       (p1_dl[8]    )
   );

   (* BEL="X11/Y2/lc0" *)
   SB_DFF  dff_3_8 (
      .C       (i_clk         ),
      .D       (p1_dl[8]    ),
      .Q       (o_data[8]   )
   );

   (* BEL="X10/Y2/lc1" *)
   SB_DFF  dff_2_9 (
      .C       (i_clk         ),
      .D       (p0_dl[10]  ),
      .Q       (p1_dl[9]    )
   );

   (* BEL="X11/Y2/lc1" *)
   SB_DFF  dff_3_9 (
      .C       (i_clk         ),
      .D       (p1_dl[9]    ),
      .Q       (o_data[9]   )
   );

   (* BEL="X10/Y2/lc2" *)
   SB_DFF  dff_2_10 (
      .C       (i_clk         ),
      .D       (p0_dl[11]  ),
      .Q       (p1_dl[10]    )
   );

   (* BEL="X11/Y2/lc2" *)
   SB_DFF  dff_3_10 (
      .C       (i_clk         ),
      .D       (p1_dl[10]    ),
      .Q       (o_data[10]   )
   );

   (* BEL="X10/Y2/lc3" *)
   SB_DFF  dff_2_11 (
      .C       (i_clk         ),
      .D       (p0_dl[12]  ),
      .Q       (p1_dl[11]    )
   );

   (* BEL="X11/Y2/lc3" *)
   SB_DFF  dff_3_11 (
      .C       (i_clk         ),
      .D       (p1_dl[11]    ),
      .Q       (o_data[11]   )
   );

   (* BEL="X10/Y2/lc4" *)
   SB_DFF  dff_2_12 (
      .C       (i_clk         ),
      .D       (p0_dl[13]  ),
      .Q       (p1_dl[12]    )
   );

   (* BEL="X11/Y2/lc4" *)
   SB_DFF  dff_3_12 (
      .C       (i_clk         ),
      .D       (p1_dl[12]    ),
      .Q       (o_data[12]   )
   );

   (* BEL="X10/Y2/lc5" *)
   SB_DFF  dff_2_13 (
      .C       (i_clk         ),
      .D       (p0_dl[14]  ),
      .Q       (p1_dl[13]    )
   );

   (* BEL="X11/Y2/lc5" *)
   SB_DFF  dff_3_13 (
      .C       (i_clk         ),
      .D       (p1_dl[13]    ),
      .Q       (o_data[13]   )
   );

   (* BEL="X10/Y2/lc6" *)
   SB_DFF  dff_2_14 (
      .C       (i_clk         ),
      .D       (p0_dl[15]  ),
      .Q       (p1_dl[14]    )
   );

   (* BEL="X11/Y2/lc6" *)
   SB_DFF  dff_3_14 (
      .C       (i_clk         ),
      .D       (p1_dl[14]    ),
      .Q       (o_data[14]   )
   );

   (* BEL="X10/Y2/lc7" *)
   SB_DFF  dff_2_15 (
      .C       (i_clk         ),
      .D       (p0_dl[16]  ),
      .Q       (p1_dl[15]    )
   );

   (* BEL="X11/Y2/lc7" *)
   SB_DFF  dff_3_15 (
      .C       (i_clk         ),
      .D       (p1_dl[15]    ),
      .Q       (o_data[15]   )
   );

   (* BEL="X10/Y3/lc0" *)
   SB_DFF  dff_2_16 (
      .C       (i_clk         ),
      .D       (p0_dl[17]  ),
      .Q       (p1_dl[16]    )
   );

   (* BEL="X11/Y3/lc0" *)
   SB_DFF  dff_3_16 (
      .C       (i_clk         ),
      .D       (p1_dl[16]    ),
      .Q       (o_data[16]   )
   );

   (* BEL="X10/Y3/lc1" *)
   SB_DFF  dff_2_17 (
      .C       (i_clk         ),
      .D       (p0_dl[18]  ),
      .Q       (p1_dl[17]    )
   );

   (* BEL="X11/Y3/lc1" *)
   SB_DFF  dff_3_17 (
      .C       (i_clk         ),
      .D       (p1_dl[17]    ),
      .Q       (o_data[17]   )
   );

   (* BEL="X10/Y3/lc2" *)
   SB_DFF  dff_2_18 (
      .C       (i_clk         ),
      .D       (p0_dl[19]  ),
      .Q       (p1_dl[18]    )
   );

   (* BEL="X11/Y3/lc2" *)
   SB_DFF  dff_3_18 (
      .C       (i_clk         ),
      .D       (p1_dl[18]    ),
      .Q       (o_data[18]   )
   );

   (* BEL="X10/Y3/lc3" *)
   SB_DFF  dff_2_19 (
      .C       (i_clk         ),
      .D       (p0_dl[20]  ),
      .Q       (p1_dl[19]    )
   );

   (* BEL="X11/Y3/lc3" *)
   SB_DFF  dff_3_19 (
      .C       (i_clk         ),
      .D       (p1_dl[19]    ),
      .Q       (o_data[19]   )
   );

   (* BEL="X10/Y3/lc4" *)
   SB_DFF  dff_2_20 (
      .C       (i_clk         ),
      .D       (p0_dl[21]  ),
      .Q       (p1_dl[20]    )
   );

   (* BEL="X11/Y3/lc4" *)
   SB_DFF  dff_3_20 (
      .C       (i_clk         ),
      .D       (p1_dl[20]    ),
      .Q       (o_data[20]   )
   );

   (* BEL="X10/Y3/lc5" *)
   SB_DFF  dff_2_21 (
      .C       (i_clk         ),
      .D       (p0_dl[22]  ),
      .Q       (p1_dl[21]    )
   );

   (* BEL="X11/Y3/lc5" *)
   SB_DFF  dff_3_21 (
      .C       (i_clk         ),
      .D       (p1_dl[21]    ),
      .Q       (o_data[21]   )
   );

   (* BEL="X10/Y3/lc6" *)
   SB_DFF  dff_2_22 (
      .C       (i_clk         ),
      .D       (p0_dl[23]  ),
      .Q       (p1_dl[22]    )
   );

   (* BEL="X11/Y3/lc6" *)
   SB_DFF  dff_3_22 (
      .C       (i_clk         ),
      .D       (p1_dl[22]    ),
      .Q       (o_data[22]   )
   );

   (* BEL="X10/Y3/lc7" *)
   SB_DFF  dff_2_23 (
      .C       (i_clk         ),
      .D       (p0_dl[24]  ),
      .Q       (p1_dl[23]    )
   );

   (* BEL="X11/Y3/lc7" *)
   SB_DFF  dff_3_23 (
      .C       (i_clk         ),
      .D       (p1_dl[23]    ),
      .Q       (o_data[23]   )
   );

   (* BEL="X10/Y4/lc0" *)
   SB_DFF  dff_2_24 (
      .C       (i_clk         ),
      .D       (p0_dl[25]  ),
      .Q       (p1_dl[24]    )
   );

   (* BEL="X11/Y4/lc0" *)
   SB_DFF  dff_3_24 (
      .C       (i_clk         ),
      .D       (p1_dl[24]    ),
      .Q       (o_data[24]   )
   );

   (* BEL="X10/Y4/lc1" *)
   SB_DFF  dff_2_25 (
      .C       (i_clk         ),
      .D       (p0_dl[26]  ),
      .Q       (p1_dl[25]    )
   );

   (* BEL="X11/Y4/lc1" *)
   SB_DFF  dff_3_25 (
      .C       (i_clk         ),
      .D       (p1_dl[25]    ),
      .Q       (o_data[25]   )
   );

   (* BEL="X10/Y4/lc2" *)
   SB_DFF  dff_2_26 (
      .C       (i_clk         ),
      .D       (p0_dl[27]  ),
      .Q       (p1_dl[26]    )
   );

   (* BEL="X11/Y4/lc2" *)
   SB_DFF  dff_3_26 (
      .C       (i_clk         ),
      .D       (p1_dl[26]    ),
      .Q       (o_data[26]   )
   );

   (* BEL="X10/Y4/lc3" *)
   SB_DFF  dff_2_27 (
      .C       (i_clk         ),
      .D       (p0_dl[28]  ),
      .Q       (p1_dl[27]    )
   );

   (* BEL="X11/Y4/lc3" *)
   SB_DFF  dff_3_27 (
      .C       (i_clk         ),
      .D       (p1_dl[27]    ),
      .Q       (o_data[27]   )
   );

   (* BEL="X10/Y4/lc4" *)
   SB_DFF  dff_2_28 (
      .C       (i_clk         ),
      .D       (p0_dl[29]  ),
      .Q       (p1_dl[28]    )
   );

   (* BEL="X11/Y4/lc4" *)
   SB_DFF  dff_3_28 (
      .C       (i_clk         ),
      .D       (p1_dl[28]    ),
      .Q       (o_data[28]   )
   );

   (* BEL="X10/Y4/lc5" *)
   SB_DFF  dff_2_29 (
      .C       (i_clk         ),
      .D       (p0_dl[30]  ),
      .Q       (p1_dl[29]    )
   );

   (* BEL="X11/Y4/lc5" *)
   SB_DFF  dff_3_29 (
      .C       (i_clk         ),
      .D       (p1_dl[29]    ),
      .Q       (o_data[29]   )
   );

   (* BEL="X10/Y4/lc6" *)
   SB_DFF  dff_2_30 (
      .C       (i_clk         ),
      .D       (p0_dl[31]  ),
      .Q       (p1_dl[30]    )
   );

   (* BEL="X11/Y4/lc6" *)
   SB_DFF  dff_3_30 (
      .C       (i_clk         ),
      .D       (p1_dl[30]    ),
      .Q       (o_data[30]   )
   );

   (* BEL="X10/Y4/lc7" *)
   SB_DFF  dff_2_31 (
      .C       (i_clk         ),
      .D       (p0_dl[32]  ),
      .Q       (p1_dl[31]    )
   );

   (* BEL="X11/Y4/lc7" *)
   SB_DFF  dff_3_31 (
      .C       (i_clk         ),
      .D       (p1_dl[31]    ),
      .Q       (o_data[31]   )
   );

   (* BEL="X10/Y5/lc0" *)
   SB_DFF  dff_2_32 (
      .C       (i_clk         ),
      .D       (p0_dl[33]  ),
      .Q       (p1_dl[32]    )
   );

   (* BEL="X11/Y5/lc0" *)
   SB_DFF  dff_3_32 (
      .C       (i_clk         ),
      .D       (p1_dl[32]    ),
      .Q       (o_data[32]   )
   );

   (* BEL="X10/Y5/lc1" *)
   SB_DFF  dff_2_33 (
      .C       (i_clk         ),
      .D       (p0_dl[34]  ),
      .Q       (p1_dl[33]    )
   );

   (* BEL="X11/Y5/lc1" *)
   SB_DFF  dff_3_33 (
      .C       (i_clk         ),
      .D       (p1_dl[33]    ),
      .Q       (o_data[33]   )
   );

   (* BEL="X10/Y5/lc2" *)
   SB_DFF  dff_2_34 (
      .C       (i_clk         ),
      .D       (p0_dl[35]  ),
      .Q       (p1_dl[34]    )
   );

   (* BEL="X11/Y5/lc2" *)
   SB_DFF  dff_3_34 (
      .C       (i_clk         ),
      .D       (p1_dl[34]    ),
      .Q       (o_data[34]   )
   );

   (* BEL="X10/Y5/lc3" *)
   SB_DFF  dff_2_35 (
      .C       (i_clk         ),
      .D       (p0_dl[36]  ),
      .Q       (p1_dl[35]    )
   );

   (* BEL="X11/Y5/lc3" *)
   SB_DFF  dff_3_35 (
      .C       (i_clk         ),
      .D       (p1_dl[35]    ),
      .Q       (o_data[35]   )
   );

   (* BEL="X10/Y5/lc4" *)
   SB_DFF  dff_2_36 (
      .C       (i_clk         ),
      .D       (p0_dl[37]  ),
      .Q       (p1_dl[36]    )
   );

   (* BEL="X11/Y5/lc4" *)
   SB_DFF  dff_3_36 (
      .C       (i_clk         ),
      .D       (p1_dl[36]    ),
      .Q       (o_data[36]   )
   );

   (* BEL="X10/Y5/lc5" *)
   SB_DFF  dff_2_37 (
      .C       (i_clk         ),
      .D       (p0_dl[38]  ),
      .Q       (p1_dl[37]    )
   );

   (* BEL="X11/Y5/lc5" *)
   SB_DFF  dff_3_37 (
      .C       (i_clk         ),
      .D       (p1_dl[37]    ),
      .Q       (o_data[37]   )
   );

   (* BEL="X10/Y5/lc6" *)
   SB_DFF  dff_2_38 (
      .C       (i_clk         ),
      .D       (p0_dl[39]  ),
      .Q       (p1_dl[38]    )
   );

   (* BEL="X11/Y5/lc6" *)
   SB_DFF  dff_3_38 (
      .C       (i_clk         ),
      .D       (p1_dl[38]    ),
      .Q       (o_data[38]   )
   );

   (* BEL="X10/Y5/lc7" *)
   SB_DFF  dff_2_39 (
      .C       (i_clk         ),
      .D       (p0_dl[40]  ),
      .Q       (p1_dl[39]    )
   );

   (* BEL="X11/Y5/lc7" *)
   SB_DFF  dff_3_39 (
      .C       (i_clk         ),
      .D       (p1_dl[39]    ),
      .Q       (o_data[39]   )
   );

   (* BEL="X10/Y6/lc0" *)
   SB_DFF  dff_2_40 (
      .C       (i_clk         ),
      .D       (p0_dl[41]  ),
      .Q       (p1_dl[40]    )
   );

   (* BEL="X11/Y6/lc0" *)
   SB_DFF  dff_3_40 (
      .C       (i_clk         ),
      .D       (p1_dl[40]    ),
      .Q       (o_data[40]   )
   );

   (* BEL="X10/Y6/lc1" *)
   SB_DFF  dff_2_41 (
      .C       (i_clk         ),
      .D       (p0_dl[42]  ),
      .Q       (p1_dl[41]    )
   );

   (* BEL="X11/Y6/lc1" *)
   SB_DFF  dff_3_41 (
      .C       (i_clk         ),
      .D       (p1_dl[41]    ),
      .Q       (o_data[41]   )
   );

   (* BEL="X10/Y6/lc2" *)
   SB_DFF  dff_2_42 (
      .C       (i_clk         ),
      .D       (p0_dl[43]  ),
      .Q       (p1_dl[42]    )
   );

   (* BEL="X11/Y6/lc2" *)
   SB_DFF  dff_3_42 (
      .C       (i_clk         ),
      .D       (p1_dl[42]    ),
      .Q       (o_data[42]   )
   );

   (* BEL="X10/Y6/lc3" *)
   SB_DFF  dff_2_43 (
      .C       (i_clk         ),
      .D       (p0_dl[44]  ),
      .Q       (p1_dl[43]    )
   );

   (* BEL="X11/Y6/lc3" *)
   SB_DFF  dff_3_43 (
      .C       (i_clk         ),
      .D       (p1_dl[43]    ),
      .Q       (o_data[43]   )
   );

   (* BEL="X10/Y6/lc4" *)
   SB_DFF  dff_2_44 (
      .C       (i_clk         ),
      .D       (p0_dl[45]  ),
      .Q       (p1_dl[44]    )
   );

   (* BEL="X11/Y6/lc4" *)
   SB_DFF  dff_3_44 (
      .C       (i_clk         ),
      .D       (p1_dl[44]    ),
      .Q       (o_data[44]   )
   );

   (* BEL="X10/Y6/lc5" *)
   SB_DFF  dff_2_45 (
      .C       (i_clk         ),
      .D       (p0_dl[46]  ),
      .Q       (p1_dl[45]    )
   );

   (* BEL="X11/Y6/lc5" *)
   SB_DFF  dff_3_45 (
      .C       (i_clk         ),
      .D       (p1_dl[45]    ),
      .Q       (o_data[45]   )
   );

   (* BEL="X10/Y6/lc6" *)
   SB_DFF  dff_2_46 (
      .C       (i_clk         ),
      .D       (p0_dl[47]  ),
      .Q       (p1_dl[46]    )
   );

   (* BEL="X11/Y6/lc6" *)
   SB_DFF  dff_3_46 (
      .C       (i_clk         ),
      .D       (p1_dl[46]    ),
      .Q       (o_data[46]   )
   );

   (* BEL="X10/Y6/lc7" *)
   SB_DFF  dff_2_47 (
      .C       (i_clk         ),
      .D       (p0_dl[48]  ),
      .Q       (p1_dl[47]    )
   );

   (* BEL="X11/Y6/lc7" *)
   SB_DFF  dff_3_47 (
      .C       (i_clk         ),
      .D       (p1_dl[47]    ),
      .Q       (o_data[47]   )
   );

   (* BEL="X10/Y7/lc0" *)
   SB_DFF  dff_2_48 (
      .C       (i_clk         ),
      .D       (p0_dl[49]  ),
      .Q       (p1_dl[48]    )
   );

   (* BEL="X11/Y7/lc0" *)
   SB_DFF  dff_3_48 (
      .C       (i_clk         ),
      .D       (p1_dl[48]    ),
      .Q       (o_data[48]   )
   );

   (* BEL="X10/Y7/lc1" *)
   SB_DFF  dff_2_49 (
      .C       (i_clk         ),
      .D       (p0_dl[50]  ),
      .Q       (p1_dl[49]    )
   );

   (* BEL="X11/Y7/lc1" *)
   SB_DFF  dff_3_49 (
      .C       (i_clk         ),
      .D       (p1_dl[49]    ),
      .Q       (o_data[49]   )
   );

   (* BEL="X10/Y7/lc2" *)
   SB_DFF  dff_2_50 (
      .C       (i_clk         ),
      .D       (p0_dl[51]  ),
      .Q       (p1_dl[50]    )
   );

   (* BEL="X11/Y7/lc2" *)
   SB_DFF  dff_3_50 (
      .C       (i_clk         ),
      .D       (p1_dl[50]    ),
      .Q       (o_data[50]   )
   );

   (* BEL="X10/Y7/lc3" *)
   SB_DFF  dff_2_51 (
      .C       (i_clk         ),
      .D       (p0_dl[52]  ),
      .Q       (p1_dl[51]    )
   );

   (* BEL="X11/Y7/lc3" *)
   SB_DFF  dff_3_51 (
      .C       (i_clk         ),
      .D       (p1_dl[51]    ),
      .Q       (o_data[51]   )
   );

   (* BEL="X10/Y7/lc4" *)
   SB_DFF  dff_2_52 (
      .C       (i_clk         ),
      .D       (p0_dl[53]  ),
      .Q       (p1_dl[52]    )
   );

   (* BEL="X11/Y7/lc4" *)
   SB_DFF  dff_3_52 (
      .C       (i_clk         ),
      .D       (p1_dl[52]    ),
      .Q       (o_data[52]   )
   );

   (* BEL="X10/Y7/lc5" *)
   SB_DFF  dff_2_53 (
      .C       (i_clk         ),
      .D       (p0_dl[54]  ),
      .Q       (p1_dl[53]    )
   );

   (* BEL="X11/Y7/lc5" *)
   SB_DFF  dff_3_53 (
      .C       (i_clk         ),
      .D       (p1_dl[53]    ),
      .Q       (o_data[53]   )
   );

   (* BEL="X10/Y7/lc6" *)
   SB_DFF  dff_2_54 (
      .C       (i_clk         ),
      .D       (p0_dl[55]  ),
      .Q       (p1_dl[54]    )
   );

   (* BEL="X11/Y7/lc6" *)
   SB_DFF  dff_3_54 (
      .C       (i_clk         ),
      .D       (p1_dl[54]    ),
      .Q       (o_data[54]   )
   );

   (* BEL="X10/Y7/lc7" *)
   SB_DFF  dff_2_55 (
      .C       (i_clk         ),
      .D       (p0_dl[56]  ),
      .Q       (p1_dl[55]    )
   );

   (* BEL="X11/Y7/lc7" *)
   SB_DFF  dff_3_55 (
      .C       (i_clk         ),
      .D       (p1_dl[55]    ),
      .Q       (o_data[55]   )
   );

   (* BEL="X10/Y8/lc0" *)
   SB_DFF  dff_2_56 (
      .C       (i_clk         ),
      .D       (p0_dl[57]  ),
      .Q       (p1_dl[56]    )
   );

   (* BEL="X11/Y8/lc0" *)
   SB_DFF  dff_3_56 (
      .C       (i_clk         ),
      .D       (p1_dl[56]    ),
      .Q       (o_data[56]   )
   );

   (* BEL="X10/Y8/lc1" *)
   SB_DFF  dff_2_57 (
      .C       (i_clk         ),
      .D       (p0_dl[58]  ),
      .Q       (p1_dl[57]    )
   );

   (* BEL="X11/Y8/lc1" *)
   SB_DFF  dff_3_57 (
      .C       (i_clk         ),
      .D       (p1_dl[57]    ),
      .Q       (o_data[57]   )
   );

   (* BEL="X10/Y8/lc2" *)
   SB_DFF  dff_2_58 (
      .C       (i_clk         ),
      .D       (p0_dl[59]  ),
      .Q       (p1_dl[58]    )
   );

   (* BEL="X11/Y8/lc2" *)
   SB_DFF  dff_3_58 (
      .C       (i_clk         ),
      .D       (p1_dl[58]    ),
      .Q       (o_data[58]   )
   );

   (* BEL="X10/Y8/lc3" *)
   SB_DFF  dff_2_59 (
      .C       (i_clk         ),
      .D       (p0_dl[60]  ),
      .Q       (p1_dl[59]    )
   );

   (* BEL="X11/Y8/lc3" *)
   SB_DFF  dff_3_59 (
      .C       (i_clk         ),
      .D       (p1_dl[59]    ),
      .Q       (o_data[59]   )
   );

   (* BEL="X10/Y8/lc4" *)
   SB_DFF  dff_2_60 (
      .C       (i_clk         ),
      .D       (p0_dl[61]  ),
      .Q       (p1_dl[60]    )
   );

   (* BEL="X11/Y8/lc4" *)
   SB_DFF  dff_3_60 (
      .C       (i_clk         ),
      .D       (p1_dl[60]    ),
      .Q       (o_data[60]   )
   );

   (* BEL="X10/Y8/lc5" *)
   SB_DFF  dff_2_61 (
      .C       (i_clk         ),
      .D       (p0_dl[62]  ),
      .Q       (p1_dl[61]    )
   );

   (* BEL="X11/Y8/lc5" *)
   SB_DFF  dff_3_61 (
      .C       (i_clk         ),
      .D       (p1_dl[61]    ),
      .Q       (o_data[61]   )
   );

   (* BEL="X10/Y8/lc6" *)
   SB_DFF  dff_2_62 (
      .C       (i_clk         ),
      .D       (p0_dl[63]  ),
      .Q       (p1_dl[62]    )
   );

   (* BEL="X11/Y8/lc6" *)
   SB_DFF  dff_3_62 (
      .C       (i_clk         ),
      .D       (p1_dl[62]    ),
      .Q       (o_data[62]   )
   );

   (* BEL="X10/Y8/lc7" *)
   SB_DFF  dff_2_63 (
      .C       (i_clk         ),
      .D       (p0_dl[64]  ),
      .Q       (p1_dl[63]    )
   );

   (* BEL="X11/Y8/lc7" *)
   SB_DFF  dff_3_63 (
      .C       (i_clk         ),
      .D       (p1_dl[63]    ),
      .Q       (o_data[63]   )
   );

   (* BEL="X10/Y9/lc0" *)
   SB_DFF  dff_2_64 (
      .C       (i_clk         ),
      .D       (p0_dl[65]  ),
      .Q       (p1_dl[64]    )
   );

   (* BEL="X11/Y9/lc0" *)
   SB_DFF  dff_3_64 (
      .C       (i_clk         ),
      .D       (p1_dl[64]    ),
      .Q       (o_data[64]   )
   );

   (* BEL="X10/Y9/lc1" *)
   SB_DFF  dff_2_65 (
      .C       (i_clk         ),
      .D       (p0_dl[66]  ),
      .Q       (p1_dl[65]    )
   );

   (* BEL="X11/Y9/lc1" *)
   SB_DFF  dff_3_65 (
      .C       (i_clk         ),
      .D       (p1_dl[65]    ),
      .Q       (o_data[65]   )
   );

   (* BEL="X10/Y9/lc2" *)
   SB_DFF  dff_2_66 (
      .C       (i_clk         ),
      .D       (p0_dl[67]  ),
      .Q       (p1_dl[66]    )
   );

   (* BEL="X11/Y9/lc2" *)
   SB_DFF  dff_3_66 (
      .C       (i_clk         ),
      .D       (p1_dl[66]    ),
      .Q       (o_data[66]   )
   );

   (* BEL="X10/Y9/lc3" *)
   SB_DFF  dff_2_67 (
      .C       (i_clk         ),
      .D       (p0_dl[68]  ),
      .Q       (p1_dl[67]    )
   );

   (* BEL="X11/Y9/lc3" *)
   SB_DFF  dff_3_67 (
      .C       (i_clk         ),
      .D       (p1_dl[67]    ),
      .Q       (o_data[67]   )
   );

   (* BEL="X10/Y9/lc4" *)
   SB_DFF  dff_2_68 (
      .C       (i_clk         ),
      .D       (p0_dl[69]  ),
      .Q       (p1_dl[68]    )
   );

   (* BEL="X11/Y9/lc4" *)
   SB_DFF  dff_3_68 (
      .C       (i_clk         ),
      .D       (p1_dl[68]    ),
      .Q       (o_data[68]   )
   );

   (* BEL="X10/Y9/lc5" *)
   SB_DFF  dff_2_69 (
      .C       (i_clk         ),
      .D       (p0_dl[70]  ),
      .Q       (p1_dl[69]    )
   );

   (* BEL="X11/Y9/lc5" *)
   SB_DFF  dff_3_69 (
      .C       (i_clk         ),
      .D       (p1_dl[69]    ),
      .Q       (o_data[69]   )
   );

   (* BEL="X10/Y9/lc6" *)
   SB_DFF  dff_2_70 (
      .C       (i_clk         ),
      .D       (p0_dl[71]  ),
      .Q       (p1_dl[70]    )
   );

   (* BEL="X11/Y9/lc6" *)
   SB_DFF  dff_3_70 (
      .C       (i_clk         ),
      .D       (p1_dl[70]    ),
      .Q       (o_data[70]   )
   );

   (* BEL="X10/Y9/lc7" *)
   SB_DFF  dff_2_71 (
      .C       (i_clk         ),
      .D       (p0_dl[72]  ),
      .Q       (p1_dl[71]    )
   );

   (* BEL="X11/Y9/lc7" *)
   SB_DFF  dff_3_71 (
      .C       (i_clk         ),
      .D       (p1_dl[71]    ),
      .Q       (o_data[71]   )
   );

   (* BEL="X10/Y10/lc0" *)
   SB_DFF  dff_2_72 (
      .C       (i_clk         ),
      .D       (p0_dl[73]  ),
      .Q       (p1_dl[72]    )
   );

   (* BEL="X11/Y10/lc0" *)
   SB_DFF  dff_3_72 (
      .C       (i_clk         ),
      .D       (p1_dl[72]    ),
      .Q       (o_data[72]   )
   );

   (* BEL="X10/Y10/lc1" *)
   SB_DFF  dff_2_73 (
      .C       (i_clk         ),
      .D       (p0_dl[74]  ),
      .Q       (p1_dl[73]    )
   );

   (* BEL="X11/Y10/lc1" *)
   SB_DFF  dff_3_73 (
      .C       (i_clk         ),
      .D       (p1_dl[73]    ),
      .Q       (o_data[73]   )
   );

   (* BEL="X10/Y10/lc2" *)
   SB_DFF  dff_2_74 (
      .C       (i_clk         ),
      .D       (p0_dl[75]  ),
      .Q       (p1_dl[74]    )
   );

   (* BEL="X11/Y10/lc2" *)
   SB_DFF  dff_3_74 (
      .C       (i_clk         ),
      .D       (p1_dl[74]    ),
      .Q       (o_data[74]   )
   );

   (* BEL="X10/Y10/lc3" *)
   SB_DFF  dff_2_75 (
      .C       (i_clk         ),
      .D       (p0_dl[76]  ),
      .Q       (p1_dl[75]    )
   );

   (* BEL="X11/Y10/lc3" *)
   SB_DFF  dff_3_75 (
      .C       (i_clk         ),
      .D       (p1_dl[75]    ),
      .Q       (o_data[75]   )
   );

   (* BEL="X10/Y10/lc4" *)
   SB_DFF  dff_2_76 (
      .C       (i_clk         ),
      .D       (p0_dl[77]  ),
      .Q       (p1_dl[76]    )
   );

   (* BEL="X11/Y10/lc4" *)
   SB_DFF  dff_3_76 (
      .C       (i_clk         ),
      .D       (p1_dl[76]    ),
      .Q       (o_data[76]   )
   );

   (* BEL="X10/Y10/lc5" *)
   SB_DFF  dff_2_77 (
      .C       (i_clk         ),
      .D       (p0_dl[78]  ),
      .Q       (p1_dl[77]    )
   );

   (* BEL="X11/Y10/lc5" *)
   SB_DFF  dff_3_77 (
      .C       (i_clk         ),
      .D       (p1_dl[77]    ),
      .Q       (o_data[77]   )
   );

   (* BEL="X10/Y10/lc6" *)
   SB_DFF  dff_2_78 (
      .C       (i_clk         ),
      .D       (p0_dl[79]  ),
      .Q       (p1_dl[78]    )
   );

   (* BEL="X11/Y10/lc6" *)
   SB_DFF  dff_3_78 (
      .C       (i_clk         ),
      .D       (p1_dl[78]    ),
      .Q       (o_data[78]   )
   );

   (* BEL="X10/Y10/lc7" *)
   SB_DFF  dff_2_79 (
      .C       (i_clk         ),
      .D       (p0_dl[80]  ),
      .Q       (p1_dl[79]    )
   );

   (* BEL="X11/Y10/lc7" *)
   SB_DFF  dff_3_79 (
      .C       (i_clk         ),
      .D       (p1_dl[79]    ),
      .Q       (o_data[79]   )
   );

   (* BEL="X10/Y11/lc0" *)
   SB_DFF  dff_2_80 (
      .C       (i_clk         ),
      .D       (p0_dl[81]  ),
      .Q       (p1_dl[80]    )
   );

   (* BEL="X11/Y11/lc0" *)
   SB_DFF  dff_3_80 (
      .C       (i_clk         ),
      .D       (p1_dl[80]    ),
      .Q       (o_data[80]   )
   );

   (* BEL="X10/Y11/lc1" *)
   SB_DFF  dff_2_81 (
      .C       (i_clk         ),
      .D       (p0_dl[82]  ),
      .Q       (p1_dl[81]    )
   );

   (* BEL="X11/Y11/lc1" *)
   SB_DFF  dff_3_81 (
      .C       (i_clk         ),
      .D       (p1_dl[81]    ),
      .Q       (o_data[81]   )
   );

   (* BEL="X10/Y11/lc2" *)
   SB_DFF  dff_2_82 (
      .C       (i_clk         ),
      .D       (p0_dl[83]  ),
      .Q       (p1_dl[82]    )
   );

   (* BEL="X11/Y11/lc2" *)
   SB_DFF  dff_3_82 (
      .C       (i_clk         ),
      .D       (p1_dl[82]    ),
      .Q       (o_data[82]   )
   );

   (* BEL="X10/Y11/lc3" *)
   SB_DFF  dff_2_83 (
      .C       (i_clk         ),
      .D       (p0_dl[84]  ),
      .Q       (p1_dl[83]    )
   );

   (* BEL="X11/Y11/lc3" *)
   SB_DFF  dff_3_83 (
      .C       (i_clk         ),
      .D       (p1_dl[83]    ),
      .Q       (o_data[83]   )
   );

   (* BEL="X10/Y11/lc4" *)
   SB_DFF  dff_2_84 (
      .C       (i_clk         ),
      .D       (p0_dl[85]  ),
      .Q       (p1_dl[84]    )
   );

   (* BEL="X11/Y11/lc4" *)
   SB_DFF  dff_3_84 (
      .C       (i_clk         ),
      .D       (p1_dl[84]    ),
      .Q       (o_data[84]   )
   );

   (* BEL="X10/Y11/lc5" *)
   SB_DFF  dff_2_85 (
      .C       (i_clk         ),
      .D       (p0_dl[86]  ),
      .Q       (p1_dl[85]    )
   );

   (* BEL="X11/Y11/lc5" *)
   SB_DFF  dff_3_85 (
      .C       (i_clk         ),
      .D       (p1_dl[85]    ),
      .Q       (o_data[85]   )
   );

   (* BEL="X10/Y11/lc6" *)
   SB_DFF  dff_2_86 (
      .C       (i_clk         ),
      .D       (p0_dl[87]  ),
      .Q       (p1_dl[86]    )
   );

   (* BEL="X11/Y11/lc6" *)
   SB_DFF  dff_3_86 (
      .C       (i_clk         ),
      .D       (p1_dl[86]    ),
      .Q       (o_data[86]   )
   );

   (* BEL="X10/Y11/lc7" *)
   SB_DFF  dff_2_87 (
      .C       (i_clk         ),
      .D       (p0_dl[88]  ),
      .Q       (p1_dl[87]    )
   );

   (* BEL="X11/Y11/lc7" *)
   SB_DFF  dff_3_87 (
      .C       (i_clk         ),
      .D       (p1_dl[87]    ),
      .Q       (o_data[87]   )
   );

   (* BEL="X10/Y12/lc0" *)
   SB_DFF  dff_2_88 (
      .C       (i_clk         ),
      .D       (p0_dl[89]  ),
      .Q       (p1_dl[88]    )
   );

   (* BEL="X11/Y12/lc0" *)
   SB_DFF  dff_3_88 (
      .C       (i_clk         ),
      .D       (p1_dl[88]    ),
      .Q       (o_data[88]   )
   );

   (* BEL="X10/Y12/lc1" *)
   SB_DFF  dff_2_89 (
      .C       (i_clk         ),
      .D       (p0_dl[90]  ),
      .Q       (p1_dl[89]    )
   );

   (* BEL="X11/Y12/lc1" *)
   SB_DFF  dff_3_89 (
      .C       (i_clk         ),
      .D       (p1_dl[89]    ),
      .Q       (o_data[89]   )
   );

   (* BEL="X10/Y12/lc2" *)
   SB_DFF  dff_2_90 (
      .C       (i_clk         ),
      .D       (p0_dl[91]  ),
      .Q       (p1_dl[90]    )
   );

   (* BEL="X11/Y12/lc2" *)
   SB_DFF  dff_3_90 (
      .C       (i_clk         ),
      .D       (p1_dl[90]    ),
      .Q       (o_data[90]   )
   );

   (* BEL="X10/Y12/lc3" *)
   SB_DFF  dff_2_91 (
      .C       (i_clk         ),
      .D       (p0_dl[92]  ),
      .Q       (p1_dl[91]    )
   );

   (* BEL="X11/Y12/lc3" *)
   SB_DFF  dff_3_91 (
      .C       (i_clk         ),
      .D       (p1_dl[91]    ),
      .Q       (o_data[91]   )
   );

   (* BEL="X10/Y12/lc4" *)
   SB_DFF  dff_2_92 (
      .C       (i_clk         ),
      .D       (p0_dl[93]  ),
      .Q       (p1_dl[92]    )
   );

   (* BEL="X11/Y12/lc4" *)
   SB_DFF  dff_3_92 (
      .C       (i_clk         ),
      .D       (p1_dl[92]    ),
      .Q       (o_data[92]   )
   );

   (* BEL="X10/Y12/lc5" *)
   SB_DFF  dff_2_93 (
      .C       (i_clk         ),
      .D       (p0_dl[94]  ),
      .Q       (p1_dl[93]    )
   );

   (* BEL="X11/Y12/lc5" *)
   SB_DFF  dff_3_93 (
      .C       (i_clk         ),
      .D       (p1_dl[93]    ),
      .Q       (o_data[93]   )
   );

   (* BEL="X10/Y12/lc6" *)
   SB_DFF  dff_2_94 (
      .C       (i_clk         ),
      .D       (p0_dl[95]  ),
      .Q       (p1_dl[94]    )
   );

   (* BEL="X11/Y12/lc6" *)
   SB_DFF  dff_3_94 (
      .C       (i_clk         ),
      .D       (p1_dl[94]    ),
      .Q       (o_data[94]   )
   );

   (* BEL="X10/Y12/lc7" *)
   SB_DFF  dff_2_95 (
      .C       (i_clk         ),
      .D       (p0_dl[96]  ),
      .Q       (p1_dl[95]    )
   );

   (* BEL="X11/Y12/lc7" *)
   SB_DFF  dff_3_95 (
      .C       (i_clk         ),
      .D       (p1_dl[95]    ),
      .Q       (o_data[95]   )
   );

   (* BEL="X10/Y13/lc0" *)
   SB_DFF  dff_2_96 (
      .C       (i_clk         ),
      .D       (p0_dl[97]  ),
      .Q       (p1_dl[96]    )
   );

   (* BEL="X11/Y13/lc0" *)
   SB_DFF  dff_3_96 (
      .C       (i_clk         ),
      .D       (p1_dl[96]    ),
      .Q       (o_data[96]   )
   );

   (* BEL="X10/Y13/lc1" *)
   SB_DFF  dff_2_97 (
      .C       (i_clk         ),
      .D       (p0_dl[98]  ),
      .Q       (p1_dl[97]    )
   );

   (* BEL="X11/Y13/lc1" *)
   SB_DFF  dff_3_97 (
      .C       (i_clk         ),
      .D       (p1_dl[97]    ),
      .Q       (o_data[97]   )
   );

   (* BEL="X10/Y13/lc2" *)
   SB_DFF  dff_2_98 (
      .C       (i_clk         ),
      .D       (p0_dl[99]  ),
      .Q       (p1_dl[98]    )
   );

   (* BEL="X11/Y13/lc2" *)
   SB_DFF  dff_3_98 (
      .C       (i_clk         ),
      .D       (p1_dl[98]    ),
      .Q       (o_data[98]   )
   );

   (* BEL="X10/Y13/lc3" *)
   SB_DFF  dff_2_99 (
      .C       (i_clk         ),
      .D       (p0_dl[100]  ),
      .Q       (p1_dl[99]    )
   );

   (* BEL="X11/Y13/lc3" *)
   SB_DFF  dff_3_99 (
      .C       (i_clk         ),
      .D       (p1_dl[99]    ),
      .Q       (o_data[99]   )
   );

   (* BEL="X10/Y13/lc4" *)
   SB_DFF  dff_2_100 (
      .C       (i_clk         ),
      .D       (p0_dl[101]  ),
      .Q       (p1_dl[100]    )
   );

   (* BEL="X11/Y13/lc4" *)
   SB_DFF  dff_3_100 (
      .C       (i_clk         ),
      .D       (p1_dl[100]    ),
      .Q       (o_data[100]   )
   );

   (* BEL="X10/Y13/lc5" *)
   SB_DFF  dff_2_101 (
      .C       (i_clk         ),
      .D       (p0_dl[102]  ),
      .Q       (p1_dl[101]    )
   );

   (* BEL="X11/Y13/lc5" *)
   SB_DFF  dff_3_101 (
      .C       (i_clk         ),
      .D       (p1_dl[101]    ),
      .Q       (o_data[101]   )
   );

   (* BEL="X10/Y13/lc6" *)
   SB_DFF  dff_2_102 (
      .C       (i_clk         ),
      .D       (p0_dl[103]  ),
      .Q       (p1_dl[102]    )
   );

   (* BEL="X11/Y13/lc6" *)
   SB_DFF  dff_3_102 (
      .C       (i_clk         ),
      .D       (p1_dl[102]    ),
      .Q       (o_data[102]   )
   );

   (* BEL="X10/Y13/lc7" *)
   SB_DFF  dff_2_103 (
      .C       (i_clk         ),
      .D       (p0_dl[104]  ),
      .Q       (p1_dl[103]    )
   );

   (* BEL="X11/Y13/lc7" *)
   SB_DFF  dff_3_103 (
      .C       (i_clk         ),
      .D       (p1_dl[103]    ),
      .Q       (o_data[103]   )
   );

   (* BEL="X10/Y14/lc0" *)
   SB_DFF  dff_2_104 (
      .C       (i_clk         ),
      .D       (p0_dl[105]  ),
      .Q       (p1_dl[104]    )
   );

   (* BEL="X11/Y14/lc0" *)
   SB_DFF  dff_3_104 (
      .C       (i_clk         ),
      .D       (p1_dl[104]    ),
      .Q       (o_data[104]   )
   );

   (* BEL="X10/Y14/lc1" *)
   SB_DFF  dff_2_105 (
      .C       (i_clk         ),
      .D       (p0_dl[106]  ),
      .Q       (p1_dl[105]    )
   );

   (* BEL="X11/Y14/lc1" *)
   SB_DFF  dff_3_105 (
      .C       (i_clk         ),
      .D       (p1_dl[105]    ),
      .Q       (o_data[105]   )
   );

   (* BEL="X10/Y14/lc2" *)
   SB_DFF  dff_2_106 (
      .C       (i_clk         ),
      .D       (p0_dl[107]  ),
      .Q       (p1_dl[106]    )
   );

   (* BEL="X11/Y14/lc2" *)
   SB_DFF  dff_3_106 (
      .C       (i_clk         ),
      .D       (p1_dl[106]    ),
      .Q       (o_data[106]   )
   );

   (* BEL="X10/Y14/lc3" *)
   SB_DFF  dff_2_107 (
      .C       (i_clk         ),
      .D       (p0_dl[108]  ),
      .Q       (p1_dl[107]    )
   );

   (* BEL="X11/Y14/lc3" *)
   SB_DFF  dff_3_107 (
      .C       (i_clk         ),
      .D       (p1_dl[107]    ),
      .Q       (o_data[107]   )
   );

   (* BEL="X10/Y14/lc4" *)
   SB_DFF  dff_2_108 (
      .C       (i_clk         ),
      .D       (p0_dl[109]  ),
      .Q       (p1_dl[108]    )
   );

   (* BEL="X11/Y14/lc4" *)
   SB_DFF  dff_3_108 (
      .C       (i_clk         ),
      .D       (p1_dl[108]    ),
      .Q       (o_data[108]   )
   );

   (* BEL="X10/Y14/lc5" *)
   SB_DFF  dff_2_109 (
      .C       (i_clk         ),
      .D       (p0_dl[110]  ),
      .Q       (p1_dl[109]    )
   );

   (* BEL="X11/Y14/lc5" *)
   SB_DFF  dff_3_109 (
      .C       (i_clk         ),
      .D       (p1_dl[109]    ),
      .Q       (o_data[109]   )
   );

   (* BEL="X10/Y14/lc6" *)
   SB_DFF  dff_2_110 (
      .C       (i_clk         ),
      .D       (p0_dl[111]  ),
      .Q       (p1_dl[110]    )
   );

   (* BEL="X11/Y14/lc6" *)
   SB_DFF  dff_3_110 (
      .C       (i_clk         ),
      .D       (p1_dl[110]    ),
      .Q       (o_data[110]   )
   );

   (* BEL="X10/Y14/lc7" *)
   SB_DFF  dff_2_111 (
      .C       (i_clk         ),
      .D       (p0_dl[112]  ),
      .Q       (p1_dl[111]    )
   );

   (* BEL="X11/Y14/lc7" *)
   SB_DFF  dff_3_111 (
      .C       (i_clk         ),
      .D       (p1_dl[111]    ),
      .Q       (o_data[111]   )
   );

   (* BEL="X10/Y15/lc0" *)
   SB_DFF  dff_2_112 (
      .C       (i_clk         ),
      .D       (p0_dl[113]  ),
      .Q       (p1_dl[112]    )
   );

   (* BEL="X11/Y15/lc0" *)
   SB_DFF  dff_3_112 (
      .C       (i_clk         ),
      .D       (p1_dl[112]    ),
      .Q       (o_data[112]   )
   );

   (* BEL="X10/Y15/lc1" *)
   SB_DFF  dff_2_113 (
      .C       (i_clk         ),
      .D       (p0_dl[114]  ),
      .Q       (p1_dl[113]    )
   );

   (* BEL="X11/Y15/lc1" *)
   SB_DFF  dff_3_113 (
      .C       (i_clk         ),
      .D       (p1_dl[113]    ),
      .Q       (o_data[113]   )
   );

   (* BEL="X10/Y15/lc2" *)
   SB_DFF  dff_2_114 (
      .C       (i_clk         ),
      .D       (p0_dl[115]  ),
      .Q       (p1_dl[114]    )
   );

   (* BEL="X11/Y15/lc2" *)
   SB_DFF  dff_3_114 (
      .C       (i_clk         ),
      .D       (p1_dl[114]    ),
      .Q       (o_data[114]   )
   );

   (* BEL="X10/Y15/lc3" *)
   SB_DFF  dff_2_115 (
      .C       (i_clk         ),
      .D       (p0_dl[116]  ),
      .Q       (p1_dl[115]    )
   );

   (* BEL="X11/Y15/lc3" *)
   SB_DFF  dff_3_115 (
      .C       (i_clk         ),
      .D       (p1_dl[115]    ),
      .Q       (o_data[115]   )
   );

   (* BEL="X10/Y15/lc4" *)
   SB_DFF  dff_2_116 (
      .C       (i_clk         ),
      .D       (p0_dl[117]  ),
      .Q       (p1_dl[116]    )
   );

   (* BEL="X11/Y15/lc4" *)
   SB_DFF  dff_3_116 (
      .C       (i_clk         ),
      .D       (p1_dl[116]    ),
      .Q       (o_data[116]   )
   );

   (* BEL="X10/Y15/lc5" *)
   SB_DFF  dff_2_117 (
      .C       (i_clk         ),
      .D       (p0_dl[118]  ),
      .Q       (p1_dl[117]    )
   );

   (* BEL="X11/Y15/lc5" *)
   SB_DFF  dff_3_117 (
      .C       (i_clk         ),
      .D       (p1_dl[117]    ),
      .Q       (o_data[117]   )
   );

   (* BEL="X10/Y15/lc6" *)
   SB_DFF  dff_2_118 (
      .C       (i_clk         ),
      .D       (p0_dl[119]  ),
      .Q       (p1_dl[118]    )
   );

   (* BEL="X11/Y15/lc6" *)
   SB_DFF  dff_3_118 (
      .C       (i_clk         ),
      .D       (p1_dl[118]    ),
      .Q       (o_data[118]   )
   );

   (* BEL="X10/Y15/lc7" *)
   SB_DFF  dff_2_119 (
      .C       (i_clk         ),
      .D       (p0_dl[120]  ),
      .Q       (p1_dl[119]    )
   );

   (* BEL="X11/Y15/lc7" *)
   SB_DFF  dff_3_119 (
      .C       (i_clk         ),
      .D       (p1_dl[119]    ),
      .Q       (o_data[119]   )
   );

   (* BEL="X10/Y16/lc0" *)
   SB_DFF  dff_2_120 (
      .C       (i_clk         ),
      .D       (p0_dl[121]  ),
      .Q       (p1_dl[120]    )
   );

   (* BEL="X11/Y16/lc0" *)
   SB_DFF  dff_3_120 (
      .C       (i_clk         ),
      .D       (p1_dl[120]    ),
      .Q       (o_data[120]   )
   );

   (* BEL="X10/Y16/lc1" *)
   SB_DFF  dff_2_121 (
      .C       (i_clk         ),
      .D       (p0_dl[122]  ),
      .Q       (p1_dl[121]    )
   );

   (* BEL="X11/Y16/lc1" *)
   SB_DFF  dff_3_121 (
      .C       (i_clk         ),
      .D       (p1_dl[121]    ),
      .Q       (o_data[121]   )
   );

   (* BEL="X10/Y16/lc2" *)
   SB_DFF  dff_2_122 (
      .C       (i_clk         ),
      .D       (p0_dl[123]  ),
      .Q       (p1_dl[122]    )
   );

   (* BEL="X11/Y16/lc2" *)
   SB_DFF  dff_3_122 (
      .C       (i_clk         ),
      .D       (p1_dl[122]    ),
      .Q       (o_data[122]   )
   );

   (* BEL="X10/Y16/lc3" *)
   SB_DFF  dff_2_123 (
      .C       (i_clk         ),
      .D       (p0_dl[124]  ),
      .Q       (p1_dl[123]    )
   );

   (* BEL="X11/Y16/lc3" *)
   SB_DFF  dff_3_123 (
      .C       (i_clk         ),
      .D       (p1_dl[123]    ),
      .Q       (o_data[123]   )
   );

   (* BEL="X10/Y16/lc4" *)
   SB_DFF  dff_2_124 (
      .C       (i_clk         ),
      .D       (p0_dl[125]  ),
      .Q       (p1_dl[124]    )
   );

   (* BEL="X11/Y16/lc4" *)
   SB_DFF  dff_3_124 (
      .C       (i_clk         ),
      .D       (p1_dl[124]    ),
      .Q       (o_data[124]   )
   );

   (* BEL="X10/Y16/lc5" *)
   SB_DFF  dff_2_125 (
      .C       (i_clk         ),
      .D       (p0_dl[126]  ),
      .Q       (p1_dl[125]    )
   );

   (* BEL="X11/Y16/lc5" *)
   SB_DFF  dff_3_125 (
      .C       (i_clk         ),
      .D       (p1_dl[125]    ),
      .Q       (o_data[125]   )
   );

   (* BEL="X10/Y16/lc6" *)
   SB_DFF  dff_2_126 (
      .C       (i_clk         ),
      .D       (p0_dl[127]  ),
      .Q       (p1_dl[126]    )
   );

   (* BEL="X11/Y16/lc6" *)
   SB_DFF  dff_3_126 (
      .C       (i_clk         ),
      .D       (p1_dl[126]    ),
      .Q       (o_data[126]   )
   );

   (* BEL="X10/Y16/lc7" *)
   SB_DFF  dff_2_127 (
      .C       (i_clk         ),
      .D       (p0_dl[128]  ),
      .Q       (p1_dl[127]    )
   );

   (* BEL="X11/Y16/lc7" *)
   SB_DFF  dff_3_127 (
      .C       (i_clk         ),
      .D       (p1_dl[127]    ),
      .Q       (o_data[127]   )
   );

   (* BEL="X10/Y17/lc0" *)
   SB_DFF  dff_2_128 (
      .C       (i_clk         ),
      .D       (p0_dl[129]  ),
      .Q       (p1_dl[128]    )
   );

   (* BEL="X11/Y17/lc0" *)
   SB_DFF  dff_3_128 (
      .C       (i_clk         ),
      .D       (p1_dl[128]    ),
      .Q       (o_data[128]   )
   );

   (* BEL="X10/Y17/lc1" *)
   SB_DFF  dff_2_129 (
      .C       (i_clk         ),
      .D       (p0_dl[130]  ),
      .Q       (p1_dl[129]    )
   );

   (* BEL="X11/Y17/lc1" *)
   SB_DFF  dff_3_129 (
      .C       (i_clk         ),
      .D       (p1_dl[129]    ),
      .Q       (o_data[129]   )
   );

   (* BEL="X10/Y17/lc2" *)
   SB_DFF  dff_2_130 (
      .C       (i_clk         ),
      .D       (p0_dl[131]  ),
      .Q       (p1_dl[130]    )
   );

   (* BEL="X11/Y17/lc2" *)
   SB_DFF  dff_3_130 (
      .C       (i_clk         ),
      .D       (p1_dl[130]    ),
      .Q       (o_data[130]   )
   );

   (* BEL="X10/Y17/lc3" *)
   SB_DFF  dff_2_131 (
      .C       (i_clk         ),
      .D       (p0_dl[132]  ),
      .Q       (p1_dl[131]    )
   );

   (* BEL="X11/Y17/lc3" *)
   SB_DFF  dff_3_131 (
      .C       (i_clk         ),
      .D       (p1_dl[131]    ),
      .Q       (o_data[131]   )
   );

   (* BEL="X10/Y17/lc4" *)
   SB_DFF  dff_2_132 (
      .C       (i_clk         ),
      .D       (p0_dl[133]  ),
      .Q       (p1_dl[132]    )
   );

   (* BEL="X11/Y17/lc4" *)
   SB_DFF  dff_3_132 (
      .C       (i_clk         ),
      .D       (p1_dl[132]    ),
      .Q       (o_data[132]   )
   );

   (* BEL="X10/Y17/lc5" *)
   SB_DFF  dff_2_133 (
      .C       (i_clk         ),
      .D       (p0_dl[134]  ),
      .Q       (p1_dl[133]    )
   );

   (* BEL="X11/Y17/lc5" *)
   SB_DFF  dff_3_133 (
      .C       (i_clk         ),
      .D       (p1_dl[133]    ),
      .Q       (o_data[133]   )
   );

   (* BEL="X10/Y17/lc6" *)
   SB_DFF  dff_2_134 (
      .C       (i_clk         ),
      .D       (p0_dl[135]  ),
      .Q       (p1_dl[134]    )
   );

   (* BEL="X11/Y17/lc6" *)
   SB_DFF  dff_3_134 (
      .C       (i_clk         ),
      .D       (p1_dl[134]    ),
      .Q       (o_data[134]   )
   );

   (* BEL="X10/Y17/lc7" *)
   SB_DFF  dff_2_135 (
      .C       (i_clk         ),
      .D       (p0_dl[136]  ),
      .Q       (p1_dl[135]    )
   );

   (* BEL="X11/Y17/lc7" *)
   SB_DFF  dff_3_135 (
      .C       (i_clk         ),
      .D       (p1_dl[135]    ),
      .Q       (o_data[135]   )
   );

   (* BEL="X10/Y18/lc0" *)
   SB_DFF  dff_2_136 (
      .C       (i_clk         ),
      .D       (p0_dl[137]  ),
      .Q       (p1_dl[136]    )
   );

   (* BEL="X11/Y18/lc0" *)
   SB_DFF  dff_3_136 (
      .C       (i_clk         ),
      .D       (p1_dl[136]    ),
      .Q       (o_data[136]   )
   );

   (* BEL="X10/Y18/lc1" *)
   SB_DFF  dff_2_137 (
      .C       (i_clk         ),
      .D       (p0_dl[138]  ),
      .Q       (p1_dl[137]    )
   );

   (* BEL="X11/Y18/lc1" *)
   SB_DFF  dff_3_137 (
      .C       (i_clk         ),
      .D       (p1_dl[137]    ),
      .Q       (o_data[137]   )
   );

   (* BEL="X10/Y18/lc2" *)
   SB_DFF  dff_2_138 (
      .C       (i_clk         ),
      .D       (p0_dl[139]  ),
      .Q       (p1_dl[138]    )
   );

   (* BEL="X11/Y18/lc2" *)
   SB_DFF  dff_3_138 (
      .C       (i_clk         ),
      .D       (p1_dl[138]    ),
      .Q       (o_data[138]   )
   );

   (* BEL="X10/Y18/lc3" *)
   SB_DFF  dff_2_139 (
      .C       (i_clk         ),
      .D       (p0_dl[140]  ),
      .Q       (p1_dl[139]    )
   );

   (* BEL="X11/Y18/lc3" *)
   SB_DFF  dff_3_139 (
      .C       (i_clk         ),
      .D       (p1_dl[139]    ),
      .Q       (o_data[139]   )
   );

   (* BEL="X10/Y18/lc4" *)
   SB_DFF  dff_2_140 (
      .C       (i_clk         ),
      .D       (p0_dl[141]  ),
      .Q       (p1_dl[140]    )
   );

   (* BEL="X11/Y18/lc4" *)
   SB_DFF  dff_3_140 (
      .C       (i_clk         ),
      .D       (p1_dl[140]    ),
      .Q       (o_data[140]   )
   );

   (* BEL="X10/Y18/lc5" *)
   SB_DFF  dff_2_141 (
      .C       (i_clk         ),
      .D       (p0_dl[142]  ),
      .Q       (p1_dl[141]    )
   );

   (* BEL="X11/Y18/lc5" *)
   SB_DFF  dff_3_141 (
      .C       (i_clk         ),
      .D       (p1_dl[141]    ),
      .Q       (o_data[141]   )
   );

   (* BEL="X10/Y18/lc6" *)
   SB_DFF  dff_2_142 (
      .C       (i_clk         ),
      .D       (p0_dl[143]  ),
      .Q       (p1_dl[142]    )
   );

   (* BEL="X11/Y18/lc6" *)
   SB_DFF  dff_3_142 (
      .C       (i_clk         ),
      .D       (p1_dl[142]    ),
      .Q       (o_data[142]   )
   );

   (* BEL="X10/Y18/lc7" *)
   SB_DFF  dff_2_143 (
      .C       (i_clk         ),
      .D       (p0_dl[144]  ),
      .Q       (p1_dl[143]    )
   );

   (* BEL="X11/Y18/lc7" *)
   SB_DFF  dff_3_143 (
      .C       (i_clk         ),
      .D       (p1_dl[143]    ),
      .Q       (o_data[143]   )
   );

   (* BEL="X10/Y19/lc0" *)
   SB_DFF  dff_2_144 (
      .C       (i_clk         ),
      .D       (p0_dl[145]  ),
      .Q       (p1_dl[144]    )
   );

   (* BEL="X11/Y19/lc0" *)
   SB_DFF  dff_3_144 (
      .C       (i_clk         ),
      .D       (p1_dl[144]    ),
      .Q       (o_data[144]   )
   );

   (* BEL="X10/Y19/lc1" *)
   SB_DFF  dff_2_145 (
      .C       (i_clk         ),
      .D       (p0_dl[146]  ),
      .Q       (p1_dl[145]    )
   );

   (* BEL="X11/Y19/lc1" *)
   SB_DFF  dff_3_145 (
      .C       (i_clk         ),
      .D       (p1_dl[145]    ),
      .Q       (o_data[145]   )
   );

   (* BEL="X10/Y19/lc2" *)
   SB_DFF  dff_2_146 (
      .C       (i_clk         ),
      .D       (p0_dl[147]  ),
      .Q       (p1_dl[146]    )
   );

   (* BEL="X11/Y19/lc2" *)
   SB_DFF  dff_3_146 (
      .C       (i_clk         ),
      .D       (p1_dl[146]    ),
      .Q       (o_data[146]   )
   );

   (* BEL="X10/Y19/lc3" *)
   SB_DFF  dff_2_147 (
      .C       (i_clk         ),
      .D       (p0_dl[148]  ),
      .Q       (p1_dl[147]    )
   );

   (* BEL="X11/Y19/lc3" *)
   SB_DFF  dff_3_147 (
      .C       (i_clk         ),
      .D       (p1_dl[147]    ),
      .Q       (o_data[147]   )
   );

   (* BEL="X10/Y19/lc4" *)
   SB_DFF  dff_2_148 (
      .C       (i_clk         ),
      .D       (p0_dl[149]  ),
      .Q       (p1_dl[148]    )
   );

   (* BEL="X11/Y19/lc4" *)
   SB_DFF  dff_3_148 (
      .C       (i_clk         ),
      .D       (p1_dl[148]    ),
      .Q       (o_data[148]   )
   );

   (* BEL="X10/Y19/lc5" *)
   SB_DFF  dff_2_149 (
      .C       (i_clk         ),
      .D       (p0_dl[150]  ),
      .Q       (p1_dl[149]    )
   );

   (* BEL="X11/Y19/lc5" *)
   SB_DFF  dff_3_149 (
      .C       (i_clk         ),
      .D       (p1_dl[149]    ),
      .Q       (o_data[149]   )
   );

   (* BEL="X10/Y19/lc6" *)
   SB_DFF  dff_2_150 (
      .C       (i_clk         ),
      .D       (p0_dl[151]  ),
      .Q       (p1_dl[150]    )
   );

   (* BEL="X11/Y19/lc6" *)
   SB_DFF  dff_3_150 (
      .C       (i_clk         ),
      .D       (p1_dl[150]    ),
      .Q       (o_data[150]   )
   );

   (* BEL="X10/Y19/lc7" *)
   SB_DFF  dff_2_151 (
      .C       (i_clk         ),
      .D       (p0_dl[152]  ),
      .Q       (p1_dl[151]    )
   );

   (* BEL="X11/Y19/lc7" *)
   SB_DFF  dff_3_151 (
      .C       (i_clk         ),
      .D       (p1_dl[151]    ),
      .Q       (o_data[151]   )
   );

   (* BEL="X10/Y20/lc0" *)
   SB_DFF  dff_2_152 (
      .C       (i_clk         ),
      .D       (p0_dl[153]  ),
      .Q       (p1_dl[152]    )
   );

   (* BEL="X11/Y20/lc0" *)
   SB_DFF  dff_3_152 (
      .C       (i_clk         ),
      .D       (p1_dl[152]    ),
      .Q       (o_data[152]   )
   );

   (* BEL="X10/Y20/lc1" *)
   SB_DFF  dff_2_153 (
      .C       (i_clk         ),
      .D       (p0_dl[154]  ),
      .Q       (p1_dl[153]    )
   );

   (* BEL="X11/Y20/lc1" *)
   SB_DFF  dff_3_153 (
      .C       (i_clk         ),
      .D       (p1_dl[153]    ),
      .Q       (o_data[153]   )
   );

   (* BEL="X10/Y20/lc2" *)
   SB_DFF  dff_2_154 (
      .C       (i_clk         ),
      .D       (p0_dl[155]  ),
      .Q       (p1_dl[154]    )
   );

   (* BEL="X11/Y20/lc2" *)
   SB_DFF  dff_3_154 (
      .C       (i_clk         ),
      .D       (p1_dl[154]    ),
      .Q       (o_data[154]   )
   );

   (* BEL="X10/Y20/lc3" *)
   SB_DFF  dff_2_155 (
      .C       (i_clk         ),
      .D       (p0_dl[156]  ),
      .Q       (p1_dl[155]    )
   );

   (* BEL="X11/Y20/lc3" *)
   SB_DFF  dff_3_155 (
      .C       (i_clk         ),
      .D       (p1_dl[155]    ),
      .Q       (o_data[155]   )
   );

   (* BEL="X10/Y20/lc4" *)
   SB_DFF  dff_2_156 (
      .C       (i_clk         ),
      .D       (p0_dl[157]  ),
      .Q       (p1_dl[156]    )
   );

   (* BEL="X11/Y20/lc4" *)
   SB_DFF  dff_3_156 (
      .C       (i_clk         ),
      .D       (p1_dl[156]    ),
      .Q       (o_data[156]   )
   );

   (* BEL="X10/Y20/lc5" *)
   SB_DFF  dff_2_157 (
      .C       (i_clk         ),
      .D       (p0_dl[158]  ),
      .Q       (p1_dl[157]    )
   );

   (* BEL="X11/Y20/lc5" *)
   SB_DFF  dff_3_157 (
      .C       (i_clk         ),
      .D       (p1_dl[157]    ),
      .Q       (o_data[157]   )
   );

   (* BEL="X10/Y20/lc6" *)
   SB_DFF  dff_2_158 (
      .C       (i_clk         ),
      .D       (p0_dl[159]  ),
      .Q       (p1_dl[158]    )
   );

   (* BEL="X11/Y20/lc6" *)
   SB_DFF  dff_3_158 (
      .C       (i_clk         ),
      .D       (p1_dl[158]    ),
      .Q       (o_data[158]   )
   );

   (* BEL="X10/Y20/lc7" *)
   SB_DFF  dff_2_159 (
      .C       (i_clk         ),
      .D       (p0_dl[160]  ),
      .Q       (p1_dl[159]    )
   );

   (* BEL="X11/Y20/lc7" *)
   SB_DFF  dff_3_159 (
      .C       (i_clk         ),
      .D       (p1_dl[159]    ),
      .Q       (o_data[159]   )
   );

   (* BEL="X10/Y21/lc0" *)
   SB_DFF  dff_2_160 (
      .C       (i_clk         ),
      .D       (p0_dl[161]  ),
      .Q       (p1_dl[160]    )
   );

   (* BEL="X11/Y21/lc0" *)
   SB_DFF  dff_3_160 (
      .C       (i_clk         ),
      .D       (p1_dl[160]    ),
      .Q       (o_data[160]   )
   );

   (* BEL="X10/Y21/lc1" *)
   SB_DFF  dff_2_161 (
      .C       (i_clk         ),
      .D       (p0_dl[162]  ),
      .Q       (p1_dl[161]    )
   );

   (* BEL="X11/Y21/lc1" *)
   SB_DFF  dff_3_161 (
      .C       (i_clk         ),
      .D       (p1_dl[161]    ),
      .Q       (o_data[161]   )
   );

   (* BEL="X10/Y21/lc2" *)
   SB_DFF  dff_2_162 (
      .C       (i_clk         ),
      .D       (p0_dl[163]  ),
      .Q       (p1_dl[162]    )
   );

   (* BEL="X11/Y21/lc2" *)
   SB_DFF  dff_3_162 (
      .C       (i_clk         ),
      .D       (p1_dl[162]    ),
      .Q       (o_data[162]   )
   );

   (* BEL="X10/Y21/lc3" *)
   SB_DFF  dff_2_163 (
      .C       (i_clk         ),
      .D       (p0_dl[164]  ),
      .Q       (p1_dl[163]    )
   );

   (* BEL="X11/Y21/lc3" *)
   SB_DFF  dff_3_163 (
      .C       (i_clk         ),
      .D       (p1_dl[163]    ),
      .Q       (o_data[163]   )
   );

   (* BEL="X10/Y21/lc4" *)
   SB_DFF  dff_2_164 (
      .C       (i_clk         ),
      .D       (p0_dl[165]  ),
      .Q       (p1_dl[164]    )
   );

   (* BEL="X11/Y21/lc4" *)
   SB_DFF  dff_3_164 (
      .C       (i_clk         ),
      .D       (p1_dl[164]    ),
      .Q       (o_data[164]   )
   );

   (* BEL="X10/Y21/lc5" *)
   SB_DFF  dff_2_165 (
      .C       (i_clk         ),
      .D       (p0_dl[166]  ),
      .Q       (p1_dl[165]    )
   );

   (* BEL="X11/Y21/lc5" *)
   SB_DFF  dff_3_165 (
      .C       (i_clk         ),
      .D       (p1_dl[165]    ),
      .Q       (o_data[165]   )
   );

   (* BEL="X10/Y21/lc6" *)
   SB_DFF  dff_2_166 (
      .C       (i_clk         ),
      .D       (p0_dl[167]  ),
      .Q       (p1_dl[166]    )
   );

   (* BEL="X11/Y21/lc6" *)
   SB_DFF  dff_3_166 (
      .C       (i_clk         ),
      .D       (p1_dl[166]    ),
      .Q       (o_data[166]   )
   );

   (* BEL="X10/Y21/lc7" *)
   SB_DFF  dff_2_167 (
      .C       (i_clk         ),
      .D       (p0_dl[168]  ),
      .Q       (p1_dl[167]    )
   );

   (* BEL="X11/Y21/lc7" *)
   SB_DFF  dff_3_167 (
      .C       (i_clk         ),
      .D       (p1_dl[167]    ),
      .Q       (o_data[167]   )
   );

   (* BEL="X10/Y22/lc0" *)
   SB_DFF  dff_2_168 (
      .C       (i_clk         ),
      .D       (p0_dl[169]  ),
      .Q       (p1_dl[168]    )
   );

   (* BEL="X11/Y22/lc0" *)
   SB_DFF  dff_3_168 (
      .C       (i_clk         ),
      .D       (p1_dl[168]    ),
      .Q       (o_data[168]   )
   );

   (* BEL="X10/Y22/lc1" *)
   SB_DFF  dff_2_169 (
      .C       (i_clk         ),
      .D       (p0_dl[170]  ),
      .Q       (p1_dl[169]    )
   );

   (* BEL="X11/Y22/lc1" *)
   SB_DFF  dff_3_169 (
      .C       (i_clk         ),
      .D       (p1_dl[169]    ),
      .Q       (o_data[169]   )
   );

   (* BEL="X10/Y22/lc2" *)
   SB_DFF  dff_2_170 (
      .C       (i_clk         ),
      .D       (p0_dl[171]  ),
      .Q       (p1_dl[170]    )
   );

   (* BEL="X11/Y22/lc2" *)
   SB_DFF  dff_3_170 (
      .C       (i_clk         ),
      .D       (p1_dl[170]    ),
      .Q       (o_data[170]   )
   );

   (* BEL="X10/Y22/lc3" *)
   SB_DFF  dff_2_171 (
      .C       (i_clk         ),
      .D       (p0_dl[172]  ),
      .Q       (p1_dl[171]    )
   );

   (* BEL="X11/Y22/lc3" *)
   SB_DFF  dff_3_171 (
      .C       (i_clk         ),
      .D       (p1_dl[171]    ),
      .Q       (o_data[171]   )
   );

   (* BEL="X10/Y22/lc4" *)
   SB_DFF  dff_2_172 (
      .C       (i_clk         ),
      .D       (p0_dl[173]  ),
      .Q       (p1_dl[172]    )
   );

   (* BEL="X11/Y22/lc4" *)
   SB_DFF  dff_3_172 (
      .C       (i_clk         ),
      .D       (p1_dl[172]    ),
      .Q       (o_data[172]   )
   );

   (* BEL="X10/Y22/lc5" *)
   SB_DFF  dff_2_173 (
      .C       (i_clk         ),
      .D       (p0_dl[174]  ),
      .Q       (p1_dl[173]    )
   );

   (* BEL="X11/Y22/lc5" *)
   SB_DFF  dff_3_173 (
      .C       (i_clk         ),
      .D       (p1_dl[173]    ),
      .Q       (o_data[173]   )
   );

   (* BEL="X10/Y22/lc6" *)
   SB_DFF  dff_2_174 (
      .C       (i_clk         ),
      .D       (p0_dl[175]  ),
      .Q       (p1_dl[174]    )
   );

   (* BEL="X11/Y22/lc6" *)
   SB_DFF  dff_3_174 (
      .C       (i_clk         ),
      .D       (p1_dl[174]    ),
      .Q       (o_data[174]   )
   );

   (* BEL="X10/Y22/lc7" *)
   SB_DFF  dff_2_175 (
      .C       (i_clk         ),
      .D       (p0_dl[176]  ),
      .Q       (p1_dl[175]    )
   );

   (* BEL="X11/Y22/lc7" *)
   SB_DFF  dff_3_175 (
      .C       (i_clk         ),
      .D       (p1_dl[175]    ),
      .Q       (o_data[175]   )
   );

   (* BEL="X10/Y23/lc0" *)
   SB_DFF  dff_2_176 (
      .C       (i_clk         ),
      .D       (p0_dl[177]  ),
      .Q       (p1_dl[176]    )
   );

   (* BEL="X11/Y23/lc0" *)
   SB_DFF  dff_3_176 (
      .C       (i_clk         ),
      .D       (p1_dl[176]    ),
      .Q       (o_data[176]   )
   );

   (* BEL="X10/Y23/lc1" *)
   SB_DFF  dff_2_177 (
      .C       (i_clk         ),
      .D       (p0_dl[178]  ),
      .Q       (p1_dl[177]    )
   );

   (* BEL="X11/Y23/lc1" *)
   SB_DFF  dff_3_177 (
      .C       (i_clk         ),
      .D       (p1_dl[177]    ),
      .Q       (o_data[177]   )
   );

   (* BEL="X10/Y23/lc2" *)
   SB_DFF  dff_2_178 (
      .C       (i_clk         ),
      .D       (p0_dl[179]  ),
      .Q       (p1_dl[178]    )
   );

   (* BEL="X11/Y23/lc2" *)
   SB_DFF  dff_3_178 (
      .C       (i_clk         ),
      .D       (p1_dl[178]    ),
      .Q       (o_data[178]   )
   );

   (* BEL="X10/Y23/lc3" *)
   SB_DFF  dff_2_179 (
      .C       (i_clk         ),
      .D       (p0_dl[180]  ),
      .Q       (p1_dl[179]    )
   );

   (* BEL="X11/Y23/lc3" *)
   SB_DFF  dff_3_179 (
      .C       (i_clk         ),
      .D       (p1_dl[179]    ),
      .Q       (o_data[179]   )
   );

   (* BEL="X10/Y23/lc4" *)
   SB_DFF  dff_2_180 (
      .C       (i_clk         ),
      .D       (p0_dl[181]  ),
      .Q       (p1_dl[180]    )
   );

   (* BEL="X11/Y23/lc4" *)
   SB_DFF  dff_3_180 (
      .C       (i_clk         ),
      .D       (p1_dl[180]    ),
      .Q       (o_data[180]   )
   );

   (* BEL="X10/Y23/lc5" *)
   SB_DFF  dff_2_181 (
      .C       (i_clk         ),
      .D       (p0_dl[182]  ),
      .Q       (p1_dl[181]    )
   );

   (* BEL="X11/Y23/lc5" *)
   SB_DFF  dff_3_181 (
      .C       (i_clk         ),
      .D       (p1_dl[181]    ),
      .Q       (o_data[181]   )
   );

   (* BEL="X10/Y23/lc6" *)
   SB_DFF  dff_2_182 (
      .C       (i_clk         ),
      .D       (p0_dl[183]  ),
      .Q       (p1_dl[182]    )
   );

   (* BEL="X11/Y23/lc6" *)
   SB_DFF  dff_3_182 (
      .C       (i_clk         ),
      .D       (p1_dl[182]    ),
      .Q       (o_data[182]   )
   );

   (* BEL="X10/Y23/lc7" *)
   SB_DFF  dff_2_183 (
      .C       (i_clk         ),
      .D       (p0_dl[184]  ),
      .Q       (p1_dl[183]    )
   );

   (* BEL="X11/Y23/lc7" *)
   SB_DFF  dff_3_183 (
      .C       (i_clk         ),
      .D       (p1_dl[183]    ),
      .Q       (o_data[183]   )
   );

   (* BEL="X10/Y24/lc0" *)
   SB_DFF  dff_2_184 (
      .C       (i_clk         ),
      .D       (p0_dl[185]  ),
      .Q       (p1_dl[184]    )
   );

   (* BEL="X11/Y24/lc0" *)
   SB_DFF  dff_3_184 (
      .C       (i_clk         ),
      .D       (p1_dl[184]    ),
      .Q       (o_data[184]   )
   );

   (* BEL="X10/Y24/lc1" *)
   SB_DFF  dff_2_185 (
      .C       (i_clk         ),
      .D       (p0_dl[186]  ),
      .Q       (p1_dl[185]    )
   );

   (* BEL="X11/Y24/lc1" *)
   SB_DFF  dff_3_185 (
      .C       (i_clk         ),
      .D       (p1_dl[185]    ),
      .Q       (o_data[185]   )
   );

   (* BEL="X10/Y24/lc2" *)
   SB_DFF  dff_2_186 (
      .C       (i_clk         ),
      .D       (p0_dl[187]  ),
      .Q       (p1_dl[186]    )
   );

   (* BEL="X11/Y24/lc2" *)
   SB_DFF  dff_3_186 (
      .C       (i_clk         ),
      .D       (p1_dl[186]    ),
      .Q       (o_data[186]   )
   );

   (* BEL="X10/Y24/lc3" *)
   SB_DFF  dff_2_187 (
      .C       (i_clk         ),
      .D       (p0_dl[188]  ),
      .Q       (p1_dl[187]    )
   );

   (* BEL="X11/Y24/lc3" *)
   SB_DFF  dff_3_187 (
      .C       (i_clk         ),
      .D       (p1_dl[187]    ),
      .Q       (o_data[187]   )
   );

   (* BEL="X10/Y24/lc4" *)
   SB_DFF  dff_2_188 (
      .C       (i_clk         ),
      .D       (p0_dl[189]  ),
      .Q       (p1_dl[188]    )
   );

   (* BEL="X11/Y24/lc4" *)
   SB_DFF  dff_3_188 (
      .C       (i_clk         ),
      .D       (p1_dl[188]    ),
      .Q       (o_data[188]   )
   );

   (* BEL="X10/Y24/lc5" *)
   SB_DFF  dff_2_189 (
      .C       (i_clk         ),
      .D       (p0_dl[190]  ),
      .Q       (p1_dl[189]    )
   );

   (* BEL="X11/Y24/lc5" *)
   SB_DFF  dff_3_189 (
      .C       (i_clk         ),
      .D       (p1_dl[189]    ),
      .Q       (o_data[189]   )
   );

   (* BEL="X10/Y24/lc6" *)
   SB_DFF  dff_2_190 (
      .C       (i_clk         ),
      .D       (p0_dl[191]  ),
      .Q       (p1_dl[190]    )
   );

   (* BEL="X11/Y24/lc6" *)
   SB_DFF  dff_3_190 (
      .C       (i_clk         ),
      .D       (p1_dl[190]    ),
      .Q       (o_data[190]   )
   );

   (* BEL="X10/Y24/lc7" *)
   SB_DFF  dff_2_191 (
      .C       (i_clk         ),
      .D       (p0_dl[192]  ),
      .Q       (p1_dl[191]    )
   );

   (* BEL="X11/Y24/lc7" *)
   SB_DFF  dff_3_191 (
      .C       (i_clk         ),
      .D       (p1_dl[191]    ),
      .Q       (o_data[191]   )
   );

   (* BEL="X10/Y25/lc0" *)
   SB_DFF  dff_2_192 (
      .C       (i_clk         ),
      .D       (p0_dl[193]  ),
      .Q       (p1_dl[192]    )
   );

   (* BEL="X11/Y25/lc0" *)
   SB_DFF  dff_3_192 (
      .C       (i_clk         ),
      .D       (p1_dl[192]    ),
      .Q       (o_data[192]   )
   );

   (* BEL="X10/Y25/lc1" *)
   SB_DFF  dff_2_193 (
      .C       (i_clk         ),
      .D       (p0_dl[194]  ),
      .Q       (p1_dl[193]    )
   );

   (* BEL="X11/Y25/lc1" *)
   SB_DFF  dff_3_193 (
      .C       (i_clk         ),
      .D       (p1_dl[193]    ),
      .Q       (o_data[193]   )
   );

   (* BEL="X10/Y25/lc2" *)
   SB_DFF  dff_2_194 (
      .C       (i_clk         ),
      .D       (p0_dl[195]  ),
      .Q       (p1_dl[194]    )
   );

   (* BEL="X11/Y25/lc2" *)
   SB_DFF  dff_3_194 (
      .C       (i_clk         ),
      .D       (p1_dl[194]    ),
      .Q       (o_data[194]   )
   );

   (* BEL="X10/Y25/lc3" *)
   SB_DFF  dff_2_195 (
      .C       (i_clk         ),
      .D       (p0_dl[196]  ),
      .Q       (p1_dl[195]    )
   );

   (* BEL="X11/Y25/lc3" *)
   SB_DFF  dff_3_195 (
      .C       (i_clk         ),
      .D       (p1_dl[195]    ),
      .Q       (o_data[195]   )
   );

   (* BEL="X10/Y25/lc4" *)
   SB_DFF  dff_2_196 (
      .C       (i_clk         ),
      .D       (p0_dl[197]  ),
      .Q       (p1_dl[196]    )
   );

   (* BEL="X11/Y25/lc4" *)
   SB_DFF  dff_3_196 (
      .C       (i_clk         ),
      .D       (p1_dl[196]    ),
      .Q       (o_data[196]   )
   );

   (* BEL="X10/Y25/lc5" *)
   SB_DFF  dff_2_197 (
      .C       (i_clk         ),
      .D       (p0_dl[198]  ),
      .Q       (p1_dl[197]    )
   );

   (* BEL="X11/Y25/lc5" *)
   SB_DFF  dff_3_197 (
      .C       (i_clk         ),
      .D       (p1_dl[197]    ),
      .Q       (o_data[197]   )
   );

   (* BEL="X10/Y25/lc6" *)
   SB_DFF  dff_2_198 (
      .C       (i_clk         ),
      .D       (p0_dl[199]  ),
      .Q       (p1_dl[198]    )
   );

   (* BEL="X11/Y25/lc6" *)
   SB_DFF  dff_3_198 (
      .C       (i_clk         ),
      .D       (p1_dl[198]    ),
      .Q       (o_data[198]   )
   );

   (* BEL="X10/Y25/lc7" *)
   SB_DFF  dff_2_199 (
      .C       (i_clk         ),
      .D       (p0_dl[200]  ),
      .Q       (p1_dl[199]    )
   );

   (* BEL="X11/Y25/lc7" *)
   SB_DFF  dff_3_199 (
      .C       (i_clk         ),
      .D       (p1_dl[199]    ),
      .Q       (o_data[199]   )
   );

   (* BEL="X10/Y26/lc0" *)
   SB_DFF  dff_2_200 (
      .C       (i_clk         ),
      .D       (p0_dl[201]  ),
      .Q       (p1_dl[200]    )
   );

   (* BEL="X11/Y26/lc0" *)
   SB_DFF  dff_3_200 (
      .C       (i_clk         ),
      .D       (p1_dl[200]    ),
      .Q       (o_data[200]   )
   );

   (* BEL="X10/Y26/lc1" *)
   SB_DFF  dff_2_201 (
      .C       (i_clk         ),
      .D       (p0_dl[202]  ),
      .Q       (p1_dl[201]    )
   );

   (* BEL="X11/Y26/lc1" *)
   SB_DFF  dff_3_201 (
      .C       (i_clk         ),
      .D       (p1_dl[201]    ),
      .Q       (o_data[201]   )
   );

   (* BEL="X10/Y26/lc2" *)
   SB_DFF  dff_2_202 (
      .C       (i_clk         ),
      .D       (p0_dl[203]  ),
      .Q       (p1_dl[202]    )
   );

   (* BEL="X11/Y26/lc2" *)
   SB_DFF  dff_3_202 (
      .C       (i_clk         ),
      .D       (p1_dl[202]    ),
      .Q       (o_data[202]   )
   );

   (* BEL="X10/Y26/lc3" *)
   SB_DFF  dff_2_203 (
      .C       (i_clk         ),
      .D       (p0_dl[204]  ),
      .Q       (p1_dl[203]    )
   );

   (* BEL="X11/Y26/lc3" *)
   SB_DFF  dff_3_203 (
      .C       (i_clk         ),
      .D       (p1_dl[203]    ),
      .Q       (o_data[203]   )
   );

   (* BEL="X10/Y26/lc4" *)
   SB_DFF  dff_2_204 (
      .C       (i_clk         ),
      .D       (p0_dl[205]  ),
      .Q       (p1_dl[204]    )
   );

   (* BEL="X11/Y26/lc4" *)
   SB_DFF  dff_3_204 (
      .C       (i_clk         ),
      .D       (p1_dl[204]    ),
      .Q       (o_data[204]   )
   );

   (* BEL="X10/Y26/lc5" *)
   SB_DFF  dff_2_205 (
      .C       (i_clk         ),
      .D       (p0_dl[206]  ),
      .Q       (p1_dl[205]    )
   );

   (* BEL="X11/Y26/lc5" *)
   SB_DFF  dff_3_205 (
      .C       (i_clk         ),
      .D       (p1_dl[205]    ),
      .Q       (o_data[205]   )
   );

   (* BEL="X10/Y26/lc6" *)
   SB_DFF  dff_2_206 (
      .C       (i_clk         ),
      .D       (p0_dl[207]  ),
      .Q       (p1_dl[206]    )
   );

   (* BEL="X11/Y26/lc6" *)
   SB_DFF  dff_3_206 (
      .C       (i_clk         ),
      .D       (p1_dl[206]    ),
      .Q       (o_data[206]   )
   );

   (* BEL="X10/Y26/lc7" *)
   SB_DFF  dff_2_207 (
      .C       (i_clk         ),
      .D       (p0_dl[208]  ),
      .Q       (p1_dl[207]    )
   );

   (* BEL="X11/Y26/lc7" *)
   SB_DFF  dff_3_207 (
      .C       (i_clk         ),
      .D       (p1_dl[207]    ),
      .Q       (o_data[207]   )
   );

   (* BEL="X10/Y27/lc0" *)
   SB_DFF  dff_2_208 (
      .C       (i_clk         ),
      .D       (p0_dl[209]  ),
      .Q       (p1_dl[208]    )
   );

   (* BEL="X11/Y27/lc0" *)
   SB_DFF  dff_3_208 (
      .C       (i_clk         ),
      .D       (p1_dl[208]    ),
      .Q       (o_data[208]   )
   );

   (* BEL="X10/Y27/lc1" *)
   SB_DFF  dff_2_209 (
      .C       (i_clk         ),
      .D       (p0_dl[210]  ),
      .Q       (p1_dl[209]    )
   );

   (* BEL="X11/Y27/lc1" *)
   SB_DFF  dff_3_209 (
      .C       (i_clk         ),
      .D       (p1_dl[209]    ),
      .Q       (o_data[209]   )
   );

   (* BEL="X10/Y27/lc2" *)
   SB_DFF  dff_2_210 (
      .C       (i_clk         ),
      .D       (p0_dl[211]  ),
      .Q       (p1_dl[210]    )
   );

   (* BEL="X11/Y27/lc2" *)
   SB_DFF  dff_3_210 (
      .C       (i_clk         ),
      .D       (p1_dl[210]    ),
      .Q       (o_data[210]   )
   );

   (* BEL="X10/Y27/lc3" *)
   SB_DFF  dff_2_211 (
      .C       (i_clk         ),
      .D       (p0_dl[212]  ),
      .Q       (p1_dl[211]    )
   );

   (* BEL="X11/Y27/lc3" *)
   SB_DFF  dff_3_211 (
      .C       (i_clk         ),
      .D       (p1_dl[211]    ),
      .Q       (o_data[211]   )
   );

   (* BEL="X10/Y27/lc4" *)
   SB_DFF  dff_2_212 (
      .C       (i_clk         ),
      .D       (p0_dl[213]  ),
      .Q       (p1_dl[212]    )
   );

   (* BEL="X11/Y27/lc4" *)
   SB_DFF  dff_3_212 (
      .C       (i_clk         ),
      .D       (p1_dl[212]    ),
      .Q       (o_data[212]   )
   );

   (* BEL="X10/Y27/lc5" *)
   SB_DFF  dff_2_213 (
      .C       (i_clk         ),
      .D       (p0_dl[214]  ),
      .Q       (p1_dl[213]    )
   );

   (* BEL="X11/Y27/lc5" *)
   SB_DFF  dff_3_213 (
      .C       (i_clk         ),
      .D       (p1_dl[213]    ),
      .Q       (o_data[213]   )
   );

   (* BEL="X10/Y27/lc6" *)
   SB_DFF  dff_2_214 (
      .C       (i_clk         ),
      .D       (p0_dl[215]  ),
      .Q       (p1_dl[214]    )
   );

   (* BEL="X11/Y27/lc6" *)
   SB_DFF  dff_3_214 (
      .C       (i_clk         ),
      .D       (p1_dl[214]    ),
      .Q       (o_data[214]   )
   );

   (* BEL="X10/Y27/lc7" *)
   SB_DFF  dff_2_215 (
      .C       (i_clk         ),
      .D       (p0_dl[216]  ),
      .Q       (p1_dl[215]    )
   );

   (* BEL="X11/Y27/lc7" *)
   SB_DFF  dff_3_215 (
      .C       (i_clk         ),
      .D       (p1_dl[215]    ),
      .Q       (o_data[215]   )
   );

   (* BEL="X10/Y28/lc0" *)
   SB_DFF  dff_2_216 (
      .C       (i_clk         ),
      .D       (p0_dl[217]  ),
      .Q       (p1_dl[216]    )
   );

   (* BEL="X11/Y28/lc0" *)
   SB_DFF  dff_3_216 (
      .C       (i_clk         ),
      .D       (p1_dl[216]    ),
      .Q       (o_data[216]   )
   );

   (* BEL="X10/Y28/lc1" *)
   SB_DFF  dff_2_217 (
      .C       (i_clk         ),
      .D       (p0_dl[218]  ),
      .Q       (p1_dl[217]    )
   );

   (* BEL="X11/Y28/lc1" *)
   SB_DFF  dff_3_217 (
      .C       (i_clk         ),
      .D       (p1_dl[217]    ),
      .Q       (o_data[217]   )
   );

   (* BEL="X10/Y28/lc2" *)
   SB_DFF  dff_2_218 (
      .C       (i_clk         ),
      .D       (p0_dl[219]  ),
      .Q       (p1_dl[218]    )
   );

   (* BEL="X11/Y28/lc2" *)
   SB_DFF  dff_3_218 (
      .C       (i_clk         ),
      .D       (p1_dl[218]    ),
      .Q       (o_data[218]   )
   );

   (* BEL="X10/Y28/lc3" *)
   SB_DFF  dff_2_219 (
      .C       (i_clk         ),
      .D       (p0_dl[220]  ),
      .Q       (p1_dl[219]    )
   );

   (* BEL="X11/Y28/lc3" *)
   SB_DFF  dff_3_219 (
      .C       (i_clk         ),
      .D       (p1_dl[219]    ),
      .Q       (o_data[219]   )
   );

   (* BEL="X10/Y28/lc4" *)
   SB_DFF  dff_2_220 (
      .C       (i_clk         ),
      .D       (p0_dl[221]  ),
      .Q       (p1_dl[220]    )
   );

   (* BEL="X11/Y28/lc4" *)
   SB_DFF  dff_3_220 (
      .C       (i_clk         ),
      .D       (p1_dl[220]    ),
      .Q       (o_data[220]   )
   );

   (* BEL="X10/Y28/lc5" *)
   SB_DFF  dff_2_221 (
      .C       (i_clk         ),
      .D       (p0_dl[222]  ),
      .Q       (p1_dl[221]    )
   );

   (* BEL="X11/Y28/lc5" *)
   SB_DFF  dff_3_221 (
      .C       (i_clk         ),
      .D       (p1_dl[221]    ),
      .Q       (o_data[221]   )
   );

   (* BEL="X10/Y28/lc6" *)
   SB_DFF  dff_2_222 (
      .C       (i_clk         ),
      .D       (p0_dl[223]  ),
      .Q       (p1_dl[222]    )
   );

   (* BEL="X11/Y28/lc6" *)
   SB_DFF  dff_3_222 (
      .C       (i_clk         ),
      .D       (p1_dl[222]    ),
      .Q       (o_data[222]   )
   );

   (* BEL="X10/Y28/lc7" *)
   SB_DFF  dff_2_223 (
      .C       (i_clk         ),
      .D       (p0_dl[224]  ),
      .Q       (p1_dl[223]    )
   );

   (* BEL="X11/Y28/lc7" *)
   SB_DFF  dff_3_223 (
      .C       (i_clk         ),
      .D       (p1_dl[223]    ),
      .Q       (o_data[223]   )
   );

   (* BEL="X10/Y29/lc0" *)
   SB_DFF  dff_2_224 (
      .C       (i_clk         ),
      .D       (p0_dl[225]  ),
      .Q       (p1_dl[224]    )
   );

   (* BEL="X11/Y29/lc0" *)
   SB_DFF  dff_3_224 (
      .C       (i_clk         ),
      .D       (p1_dl[224]    ),
      .Q       (o_data[224]   )
   );

   (* BEL="X10/Y29/lc1" *)
   SB_DFF  dff_2_225 (
      .C       (i_clk         ),
      .D       (p0_dl[226]  ),
      .Q       (p1_dl[225]    )
   );

   (* BEL="X11/Y29/lc1" *)
   SB_DFF  dff_3_225 (
      .C       (i_clk         ),
      .D       (p1_dl[225]    ),
      .Q       (o_data[225]   )
   );

   (* BEL="X10/Y29/lc2" *)
   SB_DFF  dff_2_226 (
      .C       (i_clk         ),
      .D       (p0_dl[227]  ),
      .Q       (p1_dl[226]    )
   );

   (* BEL="X11/Y29/lc2" *)
   SB_DFF  dff_3_226 (
      .C       (i_clk         ),
      .D       (p1_dl[226]    ),
      .Q       (o_data[226]   )
   );

   (* BEL="X10/Y29/lc3" *)
   SB_DFF  dff_2_227 (
      .C       (i_clk         ),
      .D       (p0_dl[228]  ),
      .Q       (p1_dl[227]    )
   );

   (* BEL="X11/Y29/lc3" *)
   SB_DFF  dff_3_227 (
      .C       (i_clk         ),
      .D       (p1_dl[227]    ),
      .Q       (o_data[227]   )
   );

   (* BEL="X10/Y29/lc4" *)
   SB_DFF  dff_2_228 (
      .C       (i_clk         ),
      .D       (p0_dl[229]  ),
      .Q       (p1_dl[228]    )
   );

   (* BEL="X11/Y29/lc4" *)
   SB_DFF  dff_3_228 (
      .C       (i_clk         ),
      .D       (p1_dl[228]    ),
      .Q       (o_data[228]   )
   );

   (* BEL="X10/Y29/lc5" *)
   SB_DFF  dff_2_229 (
      .C       (i_clk         ),
      .D       (p0_dl[230]  ),
      .Q       (p1_dl[229]    )
   );

   (* BEL="X11/Y29/lc5" *)
   SB_DFF  dff_3_229 (
      .C       (i_clk         ),
      .D       (p1_dl[229]    ),
      .Q       (o_data[229]   )
   );

   (* BEL="X10/Y29/lc6" *)
   SB_DFF  dff_2_230 (
      .C       (i_clk         ),
      .D       (p0_dl[231]  ),
      .Q       (p1_dl[230]    )
   );

   (* BEL="X11/Y29/lc6" *)
   SB_DFF  dff_3_230 (
      .C       (i_clk         ),
      .D       (p1_dl[230]    ),
      .Q       (o_data[230]   )
   );

   (* BEL="X10/Y29/lc7" *)
   SB_DFF  dff_2_231 (
      .C       (i_clk         ),
      .D       (p0_dl[232]  ),
      .Q       (p1_dl[231]    )
   );

   (* BEL="X11/Y29/lc7" *)
   SB_DFF  dff_3_231 (
      .C       (i_clk         ),
      .D       (p1_dl[231]    ),
      .Q       (o_data[231]   )
   );

   (* BEL="X10/Y30/lc0" *)
   SB_DFF  dff_2_232 (
      .C       (i_clk         ),
      .D       (p0_dl[233]  ),
      .Q       (p1_dl[232]    )
   );

   (* BEL="X11/Y30/lc0" *)
   SB_DFF  dff_3_232 (
      .C       (i_clk         ),
      .D       (p1_dl[232]    ),
      .Q       (o_data[232]   )
   );

   (* BEL="X10/Y30/lc1" *)
   SB_DFF  dff_2_233 (
      .C       (i_clk         ),
      .D       (p0_dl[234]  ),
      .Q       (p1_dl[233]    )
   );

   (* BEL="X11/Y30/lc1" *)
   SB_DFF  dff_3_233 (
      .C       (i_clk         ),
      .D       (p1_dl[233]    ),
      .Q       (o_data[233]   )
   );

   (* BEL="X10/Y30/lc2" *)
   SB_DFF  dff_2_234 (
      .C       (i_clk         ),
      .D       (p0_dl[235]  ),
      .Q       (p1_dl[234]    )
   );

   (* BEL="X11/Y30/lc2" *)
   SB_DFF  dff_3_234 (
      .C       (i_clk         ),
      .D       (p1_dl[234]    ),
      .Q       (o_data[234]   )
   );

   (* BEL="X10/Y30/lc3" *)
   SB_DFF  dff_2_235 (
      .C       (i_clk         ),
      .D       (p0_dl[236]  ),
      .Q       (p1_dl[235]    )
   );

   (* BEL="X11/Y30/lc3" *)
   SB_DFF  dff_3_235 (
      .C       (i_clk         ),
      .D       (p1_dl[235]    ),
      .Q       (o_data[235]   )
   );

   (* BEL="X10/Y30/lc4" *)
   SB_DFF  dff_2_236 (
      .C       (i_clk         ),
      .D       (p0_dl[237]  ),
      .Q       (p1_dl[236]    )
   );

   (* BEL="X11/Y30/lc4" *)
   SB_DFF  dff_3_236 (
      .C       (i_clk         ),
      .D       (p1_dl[236]    ),
      .Q       (o_data[236]   )
   );

   (* BEL="X10/Y30/lc5" *)
   SB_DFF  dff_2_237 (
      .C       (i_clk         ),
      .D       (p0_dl[238]  ),
      .Q       (p1_dl[237]    )
   );

   (* BEL="X11/Y30/lc5" *)
   SB_DFF  dff_3_237 (
      .C       (i_clk         ),
      .D       (p1_dl[237]    ),
      .Q       (o_data[237]   )
   );

   (* BEL="X10/Y30/lc6" *)
   SB_DFF  dff_2_238 (
      .C       (i_clk         ),
      .D       (p0_dl[239]  ),
      .Q       (p1_dl[238]    )
   );

   (* BEL="X11/Y30/lc6" *)
   SB_DFF  dff_3_238 (
      .C       (i_clk         ),
      .D       (p1_dl[238]    ),
      .Q       (o_data[238]   )
   );

   (* BEL="X10/Y30/lc7" *)
   SB_DFF  dff_2_239 (
      .C       (i_clk         ),
      .D       (p0_dl[240]  ),
      .Q       (p1_dl[239]    )
   );

   (* BEL="X11/Y30/lc7" *)
   SB_DFF  dff_3_239 (
      .C       (i_clk         ),
      .D       (p1_dl[239]    ),
      .Q       (o_data[239]   )
   );

   (* BEL="X10/Y31/lc0" *)
   SB_DFF  dff_2_240 (
      .C       (i_clk         ),
      .D       (p0_dl[241]  ),
      .Q       (p1_dl[240]    )
   );

   (* BEL="X11/Y31/lc0" *)
   SB_DFF  dff_3_240 (
      .C       (i_clk         ),
      .D       (p1_dl[240]    ),
      .Q       (o_data[240]   )
   );

   (* BEL="X10/Y31/lc1" *)
   SB_DFF  dff_2_241 (
      .C       (i_clk         ),
      .D       (p0_dl[242]  ),
      .Q       (p1_dl[241]    )
   );

   (* BEL="X11/Y31/lc1" *)
   SB_DFF  dff_3_241 (
      .C       (i_clk         ),
      .D       (p1_dl[241]    ),
      .Q       (o_data[241]   )
   );

   (* BEL="X10/Y31/lc2" *)
   SB_DFF  dff_2_242 (
      .C       (i_clk         ),
      .D       (p0_dl[243]  ),
      .Q       (p1_dl[242]    )
   );

   (* BEL="X11/Y31/lc2" *)
   SB_DFF  dff_3_242 (
      .C       (i_clk         ),
      .D       (p1_dl[242]    ),
      .Q       (o_data[242]   )
   );

   (* BEL="X10/Y31/lc3" *)
   SB_DFF  dff_2_243 (
      .C       (i_clk         ),
      .D       (p0_dl[244]  ),
      .Q       (p1_dl[243]    )
   );

   (* BEL="X11/Y31/lc3" *)
   SB_DFF  dff_3_243 (
      .C       (i_clk         ),
      .D       (p1_dl[243]    ),
      .Q       (o_data[243]   )
   );

   (* BEL="X10/Y31/lc4" *)
   SB_DFF  dff_2_244 (
      .C       (i_clk         ),
      .D       (p0_dl[245]  ),
      .Q       (p1_dl[244]    )
   );

   (* BEL="X11/Y31/lc4" *)
   SB_DFF  dff_3_244 (
      .C       (i_clk         ),
      .D       (p1_dl[244]    ),
      .Q       (o_data[244]   )
   );

   (* BEL="X10/Y31/lc5" *)
   SB_DFF  dff_2_245 (
      .C       (i_clk         ),
      .D       (p0_dl[246]  ),
      .Q       (p1_dl[245]    )
   );

   (* BEL="X11/Y31/lc5" *)
   SB_DFF  dff_3_245 (
      .C       (i_clk         ),
      .D       (p1_dl[245]    ),
      .Q       (o_data[245]   )
   );

   (* BEL="X10/Y31/lc6" *)
   SB_DFF  dff_2_246 (
      .C       (i_clk         ),
      .D       (p0_dl[247]  ),
      .Q       (p1_dl[246]    )
   );

   (* BEL="X11/Y31/lc6" *)
   SB_DFF  dff_3_246 (
      .C       (i_clk         ),
      .D       (p1_dl[246]    ),
      .Q       (o_data[246]   )
   );

   (* BEL="X10/Y31/lc7" *)
   SB_DFF  dff_2_247 (
      .C       (i_clk         ),
      .D       (p0_dl[248]  ),
      .Q       (p1_dl[247]    )
   );

   (* BEL="X11/Y31/lc7" *)
   SB_DFF  dff_3_247 (
      .C       (i_clk         ),
      .D       (p1_dl[247]    ),
      .Q       (o_data[247]   )
   );

   (* BEL="X10/Y32/lc0" *)
   SB_DFF  dff_2_248 (
      .C       (i_clk         ),
      .D       (p0_dl[249]  ),
      .Q       (p1_dl[248]    )
   );

   (* BEL="X11/Y32/lc0" *)
   SB_DFF  dff_3_248 (
      .C       (i_clk         ),
      .D       (p1_dl[248]    ),
      .Q       (o_data[248]   )
   );

   (* BEL="X10/Y32/lc1" *)
   SB_DFF  dff_2_249 (
      .C       (i_clk         ),
      .D       (p0_dl[250]  ),
      .Q       (p1_dl[249]    )
   );

   (* BEL="X11/Y32/lc1" *)
   SB_DFF  dff_3_249 (
      .C       (i_clk         ),
      .D       (p1_dl[249]    ),
      .Q       (o_data[249]   )
   );

   (* BEL="X10/Y32/lc2" *)
   SB_DFF  dff_2_250 (
      .C       (i_clk         ),
      .D       (p0_dl[251]  ),
      .Q       (p1_dl[250]    )
   );

   (* BEL="X11/Y32/lc2" *)
   SB_DFF  dff_3_250 (
      .C       (i_clk         ),
      .D       (p1_dl[250]    ),
      .Q       (o_data[250]   )
   );

   (* BEL="X10/Y32/lc3" *)
   SB_DFF  dff_2_251 (
      .C       (i_clk         ),
      .D       (p0_dl[252]  ),
      .Q       (p1_dl[251]    )
   );

   (* BEL="X11/Y32/lc3" *)
   SB_DFF  dff_3_251 (
      .C       (i_clk         ),
      .D       (p1_dl[251]    ),
      .Q       (o_data[251]   )
   );

   (* BEL="X10/Y32/lc4" *)
   SB_DFF  dff_2_252 (
      .C       (i_clk         ),
      .D       (p0_dl[253]  ),
      .Q       (p1_dl[252]    )
   );

   (* BEL="X11/Y32/lc4" *)
   SB_DFF  dff_3_252 (
      .C       (i_clk         ),
      .D       (p1_dl[252]    ),
      .Q       (o_data[252]   )
   );

   (* BEL="X10/Y32/lc5" *)
   SB_DFF  dff_2_253 (
      .C       (i_clk         ),
      .D       (p0_dl[254]  ),
      .Q       (p1_dl[253]    )
   );

   (* BEL="X11/Y32/lc5" *)
   SB_DFF  dff_3_253 (
      .C       (i_clk         ),
      .D       (p1_dl[253]    ),
      .Q       (o_data[253]   )
   );

   (* BEL="X10/Y32/lc6" *)
   SB_DFF  dff_2_254 (
      .C       (i_clk         ),
      .D       (p0_dl[255]  ),
      .Q       (p1_dl[254]    )
   );

   (* BEL="X11/Y32/lc6" *)
   SB_DFF  dff_3_254 (
      .C       (i_clk         ),
      .D       (p1_dl[254]    ),
      .Q       (o_data[254]   )
   );

   (* BEL="X10/Y32/lc7" *)
   SB_DFF  dff_2_255 (
      .C       (i_clk         ),
      .D       (p0_dl[256]  ),
      .Q       (p1_dl[255]    )
   );

   (* BEL="X11/Y32/lc7" *)
   SB_DFF  dff_3_255 (
      .C       (i_clk         ),
      .D       (p1_dl[255]    ),
      .Q       (o_data[255]   )
   );

endmodule

