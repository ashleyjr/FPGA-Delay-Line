module x_delay_line_128 (
   input    logic                         i_clk,
   input    logic                         i_dl,
   output   logic [128-1:0]          o_data
);

logic [128:0]   p0_dl;
logic [128-1:0] p1_dl;
logic [128-1:0] p2_dl;

assign p0_dl[0] = i_dl;

   (* BEL="X12/Y1/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut0 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[0]    ),
      .O       (p0_dl[1]  )
   );

   (* BEL="X12/Y1/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut1 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[1]    ),
      .O       (p0_dl[2]  )
   );

   (* BEL="X12/Y1/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut2 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[2]    ),
      .O       (p0_dl[3]  )
   );

   (* BEL="X12/Y1/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut3 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[3]    ),
      .O       (p0_dl[4]  )
   );

   (* BEL="X12/Y1/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut4 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[4]    ),
      .O       (p0_dl[5]  )
   );

   (* BEL="X12/Y1/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut5 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[5]    ),
      .O       (p0_dl[6]  )
   );

   (* BEL="X12/Y1/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut6 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[6]    ),
      .O       (p0_dl[7]  )
   );

   (* BEL="X12/Y1/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut7 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[7]    ),
      .O       (p0_dl[8]  )
   );

   (* BEL="X12/Y2/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut8 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[8]    ),
      .O       (p0_dl[9]  )
   );

   (* BEL="X12/Y2/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut9 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[9]    ),
      .O       (p0_dl[10]  )
   );

   (* BEL="X12/Y2/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut10 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[10]    ),
      .O       (p0_dl[11]  )
   );

   (* BEL="X12/Y2/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut11 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[11]    ),
      .O       (p0_dl[12]  )
   );

   (* BEL="X12/Y2/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut12 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[12]    ),
      .O       (p0_dl[13]  )
   );

   (* BEL="X12/Y2/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut13 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[13]    ),
      .O       (p0_dl[14]  )
   );

   (* BEL="X12/Y2/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut14 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[14]    ),
      .O       (p0_dl[15]  )
   );

   (* BEL="X12/Y2/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut15 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[15]    ),
      .O       (p0_dl[16]  )
   );

   (* BEL="X12/Y3/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut16 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[16]    ),
      .O       (p0_dl[17]  )
   );

   (* BEL="X12/Y3/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut17 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[17]    ),
      .O       (p0_dl[18]  )
   );

   (* BEL="X12/Y3/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut18 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[18]    ),
      .O       (p0_dl[19]  )
   );

   (* BEL="X12/Y3/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut19 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[19]    ),
      .O       (p0_dl[20]  )
   );

   (* BEL="X12/Y3/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut20 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[20]    ),
      .O       (p0_dl[21]  )
   );

   (* BEL="X12/Y3/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut21 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[21]    ),
      .O       (p0_dl[22]  )
   );

   (* BEL="X12/Y3/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut22 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[22]    ),
      .O       (p0_dl[23]  )
   );

   (* BEL="X12/Y3/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut23 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[23]    ),
      .O       (p0_dl[24]  )
   );

   (* BEL="X12/Y4/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut24 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[24]    ),
      .O       (p0_dl[25]  )
   );

   (* BEL="X12/Y4/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut25 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[25]    ),
      .O       (p0_dl[26]  )
   );

   (* BEL="X12/Y4/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut26 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[26]    ),
      .O       (p0_dl[27]  )
   );

   (* BEL="X12/Y4/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut27 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[27]    ),
      .O       (p0_dl[28]  )
   );

   (* BEL="X12/Y4/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut28 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[28]    ),
      .O       (p0_dl[29]  )
   );

   (* BEL="X12/Y4/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut29 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[29]    ),
      .O       (p0_dl[30]  )
   );

   (* BEL="X12/Y4/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut30 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[30]    ),
      .O       (p0_dl[31]  )
   );

   (* BEL="X12/Y4/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut31 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[31]    ),
      .O       (p0_dl[32]  )
   );

   (* BEL="X12/Y5/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut32 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[32]    ),
      .O       (p0_dl[33]  )
   );

   (* BEL="X12/Y5/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut33 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[33]    ),
      .O       (p0_dl[34]  )
   );

   (* BEL="X12/Y5/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut34 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[34]    ),
      .O       (p0_dl[35]  )
   );

   (* BEL="X12/Y5/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut35 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[35]    ),
      .O       (p0_dl[36]  )
   );

   (* BEL="X12/Y5/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut36 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[36]    ),
      .O       (p0_dl[37]  )
   );

   (* BEL="X12/Y5/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut37 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[37]    ),
      .O       (p0_dl[38]  )
   );

   (* BEL="X12/Y5/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut38 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[38]    ),
      .O       (p0_dl[39]  )
   );

   (* BEL="X12/Y5/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut39 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[39]    ),
      .O       (p0_dl[40]  )
   );

   (* BEL="X12/Y6/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut40 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[40]    ),
      .O       (p0_dl[41]  )
   );

   (* BEL="X12/Y6/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut41 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[41]    ),
      .O       (p0_dl[42]  )
   );

   (* BEL="X12/Y6/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut42 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[42]    ),
      .O       (p0_dl[43]  )
   );

   (* BEL="X12/Y6/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut43 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[43]    ),
      .O       (p0_dl[44]  )
   );

   (* BEL="X12/Y6/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut44 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[44]    ),
      .O       (p0_dl[45]  )
   );

   (* BEL="X12/Y6/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut45 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[45]    ),
      .O       (p0_dl[46]  )
   );

   (* BEL="X12/Y6/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut46 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[46]    ),
      .O       (p0_dl[47]  )
   );

   (* BEL="X12/Y6/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut47 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[47]    ),
      .O       (p0_dl[48]  )
   );

   (* BEL="X12/Y7/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut48 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[48]    ),
      .O       (p0_dl[49]  )
   );

   (* BEL="X12/Y7/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut49 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[49]    ),
      .O       (p0_dl[50]  )
   );

   (* BEL="X12/Y7/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut50 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[50]    ),
      .O       (p0_dl[51]  )
   );

   (* BEL="X12/Y7/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut51 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[51]    ),
      .O       (p0_dl[52]  )
   );

   (* BEL="X12/Y7/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut52 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[52]    ),
      .O       (p0_dl[53]  )
   );

   (* BEL="X12/Y7/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut53 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[53]    ),
      .O       (p0_dl[54]  )
   );

   (* BEL="X12/Y7/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut54 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[54]    ),
      .O       (p0_dl[55]  )
   );

   (* BEL="X12/Y7/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut55 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[55]    ),
      .O       (p0_dl[56]  )
   );

   (* BEL="X12/Y8/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut56 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[56]    ),
      .O       (p0_dl[57]  )
   );

   (* BEL="X12/Y8/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut57 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[57]    ),
      .O       (p0_dl[58]  )
   );

   (* BEL="X12/Y8/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut58 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[58]    ),
      .O       (p0_dl[59]  )
   );

   (* BEL="X12/Y8/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut59 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[59]    ),
      .O       (p0_dl[60]  )
   );

   (* BEL="X12/Y8/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut60 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[60]    ),
      .O       (p0_dl[61]  )
   );

   (* BEL="X12/Y8/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut61 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[61]    ),
      .O       (p0_dl[62]  )
   );

   (* BEL="X12/Y8/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut62 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[62]    ),
      .O       (p0_dl[63]  )
   );

   (* BEL="X12/Y8/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut63 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[63]    ),
      .O       (p0_dl[64]  )
   );

   (* BEL="X12/Y9/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut64 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[64]    ),
      .O       (p0_dl[65]  )
   );

   (* BEL="X12/Y9/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut65 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[65]    ),
      .O       (p0_dl[66]  )
   );

   (* BEL="X12/Y9/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut66 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[66]    ),
      .O       (p0_dl[67]  )
   );

   (* BEL="X12/Y9/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut67 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[67]    ),
      .O       (p0_dl[68]  )
   );

   (* BEL="X12/Y9/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut68 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[68]    ),
      .O       (p0_dl[69]  )
   );

   (* BEL="X12/Y9/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut69 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[69]    ),
      .O       (p0_dl[70]  )
   );

   (* BEL="X12/Y9/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut70 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[70]    ),
      .O       (p0_dl[71]  )
   );

   (* BEL="X12/Y9/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut71 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[71]    ),
      .O       (p0_dl[72]  )
   );

   (* BEL="X12/Y10/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut72 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[72]    ),
      .O       (p0_dl[73]  )
   );

   (* BEL="X12/Y10/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut73 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[73]    ),
      .O       (p0_dl[74]  )
   );

   (* BEL="X12/Y10/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut74 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[74]    ),
      .O       (p0_dl[75]  )
   );

   (* BEL="X12/Y10/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut75 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[75]    ),
      .O       (p0_dl[76]  )
   );

   (* BEL="X12/Y10/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut76 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[76]    ),
      .O       (p0_dl[77]  )
   );

   (* BEL="X12/Y10/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut77 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[77]    ),
      .O       (p0_dl[78]  )
   );

   (* BEL="X12/Y10/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut78 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[78]    ),
      .O       (p0_dl[79]  )
   );

   (* BEL="X12/Y10/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut79 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[79]    ),
      .O       (p0_dl[80]  )
   );

   (* BEL="X12/Y11/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut80 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[80]    ),
      .O       (p0_dl[81]  )
   );

   (* BEL="X12/Y11/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut81 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[81]    ),
      .O       (p0_dl[82]  )
   );

   (* BEL="X12/Y11/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut82 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[82]    ),
      .O       (p0_dl[83]  )
   );

   (* BEL="X12/Y11/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut83 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[83]    ),
      .O       (p0_dl[84]  )
   );

   (* BEL="X12/Y11/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut84 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[84]    ),
      .O       (p0_dl[85]  )
   );

   (* BEL="X12/Y11/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut85 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[85]    ),
      .O       (p0_dl[86]  )
   );

   (* BEL="X12/Y11/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut86 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[86]    ),
      .O       (p0_dl[87]  )
   );

   (* BEL="X12/Y11/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut87 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[87]    ),
      .O       (p0_dl[88]  )
   );

   (* BEL="X12/Y12/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut88 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[88]    ),
      .O       (p0_dl[89]  )
   );

   (* BEL="X12/Y12/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut89 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[89]    ),
      .O       (p0_dl[90]  )
   );

   (* BEL="X12/Y12/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut90 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[90]    ),
      .O       (p0_dl[91]  )
   );

   (* BEL="X12/Y12/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut91 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[91]    ),
      .O       (p0_dl[92]  )
   );

   (* BEL="X12/Y12/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut92 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[92]    ),
      .O       (p0_dl[93]  )
   );

   (* BEL="X12/Y12/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut93 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[93]    ),
      .O       (p0_dl[94]  )
   );

   (* BEL="X12/Y12/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut94 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[94]    ),
      .O       (p0_dl[95]  )
   );

   (* BEL="X12/Y12/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut95 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[95]    ),
      .O       (p0_dl[96]  )
   );

   (* BEL="X12/Y13/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut96 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[96]    ),
      .O       (p0_dl[97]  )
   );

   (* BEL="X12/Y13/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut97 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[97]    ),
      .O       (p0_dl[98]  )
   );

   (* BEL="X12/Y13/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut98 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[98]    ),
      .O       (p0_dl[99]  )
   );

   (* BEL="X12/Y13/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut99 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[99]    ),
      .O       (p0_dl[100]  )
   );

   (* BEL="X12/Y13/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut100 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[100]    ),
      .O       (p0_dl[101]  )
   );

   (* BEL="X12/Y13/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut101 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[101]    ),
      .O       (p0_dl[102]  )
   );

   (* BEL="X12/Y13/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut102 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[102]    ),
      .O       (p0_dl[103]  )
   );

   (* BEL="X12/Y13/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut103 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[103]    ),
      .O       (p0_dl[104]  )
   );

   (* BEL="X12/Y14/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut104 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[104]    ),
      .O       (p0_dl[105]  )
   );

   (* BEL="X12/Y14/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut105 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[105]    ),
      .O       (p0_dl[106]  )
   );

   (* BEL="X12/Y14/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut106 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[106]    ),
      .O       (p0_dl[107]  )
   );

   (* BEL="X12/Y14/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut107 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[107]    ),
      .O       (p0_dl[108]  )
   );

   (* BEL="X12/Y14/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut108 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[108]    ),
      .O       (p0_dl[109]  )
   );

   (* BEL="X12/Y14/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut109 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[109]    ),
      .O       (p0_dl[110]  )
   );

   (* BEL="X12/Y14/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut110 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[110]    ),
      .O       (p0_dl[111]  )
   );

   (* BEL="X12/Y14/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut111 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[111]    ),
      .O       (p0_dl[112]  )
   );

   (* BEL="X12/Y15/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut112 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[112]    ),
      .O       (p0_dl[113]  )
   );

   (* BEL="X12/Y15/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut113 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[113]    ),
      .O       (p0_dl[114]  )
   );

   (* BEL="X12/Y15/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut114 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[114]    ),
      .O       (p0_dl[115]  )
   );

   (* BEL="X12/Y15/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut115 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[115]    ),
      .O       (p0_dl[116]  )
   );

   (* BEL="X12/Y15/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut116 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[116]    ),
      .O       (p0_dl[117]  )
   );

   (* BEL="X12/Y15/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut117 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[117]    ),
      .O       (p0_dl[118]  )
   );

   (* BEL="X12/Y15/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut118 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[118]    ),
      .O       (p0_dl[119]  )
   );

   (* BEL="X12/Y15/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut119 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[119]    ),
      .O       (p0_dl[120]  )
   );

   (* BEL="X12/Y16/lc0" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut120 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[120]    ),
      .O       (p0_dl[121]  )
   );

   (* BEL="X12/Y16/lc1" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut121 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[121]    ),
      .O       (p0_dl[122]  )
   );

   (* BEL="X12/Y16/lc2" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut122 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[122]    ),
      .O       (p0_dl[123]  )
   );

   (* BEL="X12/Y16/lc3" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut123 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[123]    ),
      .O       (p0_dl[124]  )
   );

   (* BEL="X12/Y16/lc4" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut124 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[124]    ),
      .O       (p0_dl[125]  )
   );

   (* BEL="X12/Y16/lc5" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut125 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[125]    ),
      .O       (p0_dl[126]  )
   );

   (* BEL="X12/Y16/lc6" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut126 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[126]    ),
      .O       (p0_dl[127]  )
   );

   (* BEL="X12/Y16/lc7" *)
   SB_LUT4 #(
      .LUT_INIT(16'h0002      )
   ) lut127 (
      .I3      (1'b0          ),
      .I2      (1'b0          ),
      .I1      (1'b0          ),
      .I0      (p0_dl[127]    ),
      .O       (p0_dl[128]  )
   );


   (* BEL="X13/Y1/lc0" *)
   SB_DFF  dff_2_0 (
      .C       (i_clk         ),
      .D       (p0_dl[1]  ),
      .Q       (p1_dl[0]    )
   );

   (* BEL="X14/Y1/lc0" *)
   SB_DFF  dff_3_0 (
      .C       (i_clk         ),
      .D       (p1_dl[0]    ),
      .Q       (o_data[0]   )
   );

   (* BEL="X13/Y1/lc1" *)
   SB_DFF  dff_2_1 (
      .C       (i_clk         ),
      .D       (p0_dl[2]  ),
      .Q       (p1_dl[1]    )
   );

   (* BEL="X14/Y1/lc1" *)
   SB_DFF  dff_3_1 (
      .C       (i_clk         ),
      .D       (p1_dl[1]    ),
      .Q       (o_data[1]   )
   );

   (* BEL="X13/Y1/lc2" *)
   SB_DFF  dff_2_2 (
      .C       (i_clk         ),
      .D       (p0_dl[3]  ),
      .Q       (p1_dl[2]    )
   );

   (* BEL="X14/Y1/lc2" *)
   SB_DFF  dff_3_2 (
      .C       (i_clk         ),
      .D       (p1_dl[2]    ),
      .Q       (o_data[2]   )
   );

   (* BEL="X13/Y1/lc3" *)
   SB_DFF  dff_2_3 (
      .C       (i_clk         ),
      .D       (p0_dl[4]  ),
      .Q       (p1_dl[3]    )
   );

   (* BEL="X14/Y1/lc3" *)
   SB_DFF  dff_3_3 (
      .C       (i_clk         ),
      .D       (p1_dl[3]    ),
      .Q       (o_data[3]   )
   );

   (* BEL="X13/Y1/lc4" *)
   SB_DFF  dff_2_4 (
      .C       (i_clk         ),
      .D       (p0_dl[5]  ),
      .Q       (p1_dl[4]    )
   );

   (* BEL="X14/Y1/lc4" *)
   SB_DFF  dff_3_4 (
      .C       (i_clk         ),
      .D       (p1_dl[4]    ),
      .Q       (o_data[4]   )
   );

   (* BEL="X13/Y1/lc5" *)
   SB_DFF  dff_2_5 (
      .C       (i_clk         ),
      .D       (p0_dl[6]  ),
      .Q       (p1_dl[5]    )
   );

   (* BEL="X14/Y1/lc5" *)
   SB_DFF  dff_3_5 (
      .C       (i_clk         ),
      .D       (p1_dl[5]    ),
      .Q       (o_data[5]   )
   );

   (* BEL="X13/Y1/lc6" *)
   SB_DFF  dff_2_6 (
      .C       (i_clk         ),
      .D       (p0_dl[7]  ),
      .Q       (p1_dl[6]    )
   );

   (* BEL="X14/Y1/lc6" *)
   SB_DFF  dff_3_6 (
      .C       (i_clk         ),
      .D       (p1_dl[6]    ),
      .Q       (o_data[6]   )
   );

   (* BEL="X13/Y1/lc7" *)
   SB_DFF  dff_2_7 (
      .C       (i_clk         ),
      .D       (p0_dl[8]  ),
      .Q       (p1_dl[7]    )
   );

   (* BEL="X14/Y1/lc7" *)
   SB_DFF  dff_3_7 (
      .C       (i_clk         ),
      .D       (p1_dl[7]    ),
      .Q       (o_data[7]   )
   );

   (* BEL="X13/Y2/lc0" *)
   SB_DFF  dff_2_8 (
      .C       (i_clk         ),
      .D       (p0_dl[9]  ),
      .Q       (p1_dl[8]    )
   );

   (* BEL="X14/Y2/lc0" *)
   SB_DFF  dff_3_8 (
      .C       (i_clk         ),
      .D       (p1_dl[8]    ),
      .Q       (o_data[8]   )
   );

   (* BEL="X13/Y2/lc1" *)
   SB_DFF  dff_2_9 (
      .C       (i_clk         ),
      .D       (p0_dl[10]  ),
      .Q       (p1_dl[9]    )
   );

   (* BEL="X14/Y2/lc1" *)
   SB_DFF  dff_3_9 (
      .C       (i_clk         ),
      .D       (p1_dl[9]    ),
      .Q       (o_data[9]   )
   );

   (* BEL="X13/Y2/lc2" *)
   SB_DFF  dff_2_10 (
      .C       (i_clk         ),
      .D       (p0_dl[11]  ),
      .Q       (p1_dl[10]    )
   );

   (* BEL="X14/Y2/lc2" *)
   SB_DFF  dff_3_10 (
      .C       (i_clk         ),
      .D       (p1_dl[10]    ),
      .Q       (o_data[10]   )
   );

   (* BEL="X13/Y2/lc3" *)
   SB_DFF  dff_2_11 (
      .C       (i_clk         ),
      .D       (p0_dl[12]  ),
      .Q       (p1_dl[11]    )
   );

   (* BEL="X14/Y2/lc3" *)
   SB_DFF  dff_3_11 (
      .C       (i_clk         ),
      .D       (p1_dl[11]    ),
      .Q       (o_data[11]   )
   );

   (* BEL="X13/Y2/lc4" *)
   SB_DFF  dff_2_12 (
      .C       (i_clk         ),
      .D       (p0_dl[13]  ),
      .Q       (p1_dl[12]    )
   );

   (* BEL="X14/Y2/lc4" *)
   SB_DFF  dff_3_12 (
      .C       (i_clk         ),
      .D       (p1_dl[12]    ),
      .Q       (o_data[12]   )
   );

   (* BEL="X13/Y2/lc5" *)
   SB_DFF  dff_2_13 (
      .C       (i_clk         ),
      .D       (p0_dl[14]  ),
      .Q       (p1_dl[13]    )
   );

   (* BEL="X14/Y2/lc5" *)
   SB_DFF  dff_3_13 (
      .C       (i_clk         ),
      .D       (p1_dl[13]    ),
      .Q       (o_data[13]   )
   );

   (* BEL="X13/Y2/lc6" *)
   SB_DFF  dff_2_14 (
      .C       (i_clk         ),
      .D       (p0_dl[15]  ),
      .Q       (p1_dl[14]    )
   );

   (* BEL="X14/Y2/lc6" *)
   SB_DFF  dff_3_14 (
      .C       (i_clk         ),
      .D       (p1_dl[14]    ),
      .Q       (o_data[14]   )
   );

   (* BEL="X13/Y2/lc7" *)
   SB_DFF  dff_2_15 (
      .C       (i_clk         ),
      .D       (p0_dl[16]  ),
      .Q       (p1_dl[15]    )
   );

   (* BEL="X14/Y2/lc7" *)
   SB_DFF  dff_3_15 (
      .C       (i_clk         ),
      .D       (p1_dl[15]    ),
      .Q       (o_data[15]   )
   );

   (* BEL="X13/Y3/lc0" *)
   SB_DFF  dff_2_16 (
      .C       (i_clk         ),
      .D       (p0_dl[17]  ),
      .Q       (p1_dl[16]    )
   );

   (* BEL="X14/Y3/lc0" *)
   SB_DFF  dff_3_16 (
      .C       (i_clk         ),
      .D       (p1_dl[16]    ),
      .Q       (o_data[16]   )
   );

   (* BEL="X13/Y3/lc1" *)
   SB_DFF  dff_2_17 (
      .C       (i_clk         ),
      .D       (p0_dl[18]  ),
      .Q       (p1_dl[17]    )
   );

   (* BEL="X14/Y3/lc1" *)
   SB_DFF  dff_3_17 (
      .C       (i_clk         ),
      .D       (p1_dl[17]    ),
      .Q       (o_data[17]   )
   );

   (* BEL="X13/Y3/lc2" *)
   SB_DFF  dff_2_18 (
      .C       (i_clk         ),
      .D       (p0_dl[19]  ),
      .Q       (p1_dl[18]    )
   );

   (* BEL="X14/Y3/lc2" *)
   SB_DFF  dff_3_18 (
      .C       (i_clk         ),
      .D       (p1_dl[18]    ),
      .Q       (o_data[18]   )
   );

   (* BEL="X13/Y3/lc3" *)
   SB_DFF  dff_2_19 (
      .C       (i_clk         ),
      .D       (p0_dl[20]  ),
      .Q       (p1_dl[19]    )
   );

   (* BEL="X14/Y3/lc3" *)
   SB_DFF  dff_3_19 (
      .C       (i_clk         ),
      .D       (p1_dl[19]    ),
      .Q       (o_data[19]   )
   );

   (* BEL="X13/Y3/lc4" *)
   SB_DFF  dff_2_20 (
      .C       (i_clk         ),
      .D       (p0_dl[21]  ),
      .Q       (p1_dl[20]    )
   );

   (* BEL="X14/Y3/lc4" *)
   SB_DFF  dff_3_20 (
      .C       (i_clk         ),
      .D       (p1_dl[20]    ),
      .Q       (o_data[20]   )
   );

   (* BEL="X13/Y3/lc5" *)
   SB_DFF  dff_2_21 (
      .C       (i_clk         ),
      .D       (p0_dl[22]  ),
      .Q       (p1_dl[21]    )
   );

   (* BEL="X14/Y3/lc5" *)
   SB_DFF  dff_3_21 (
      .C       (i_clk         ),
      .D       (p1_dl[21]    ),
      .Q       (o_data[21]   )
   );

   (* BEL="X13/Y3/lc6" *)
   SB_DFF  dff_2_22 (
      .C       (i_clk         ),
      .D       (p0_dl[23]  ),
      .Q       (p1_dl[22]    )
   );

   (* BEL="X14/Y3/lc6" *)
   SB_DFF  dff_3_22 (
      .C       (i_clk         ),
      .D       (p1_dl[22]    ),
      .Q       (o_data[22]   )
   );

   (* BEL="X13/Y3/lc7" *)
   SB_DFF  dff_2_23 (
      .C       (i_clk         ),
      .D       (p0_dl[24]  ),
      .Q       (p1_dl[23]    )
   );

   (* BEL="X14/Y3/lc7" *)
   SB_DFF  dff_3_23 (
      .C       (i_clk         ),
      .D       (p1_dl[23]    ),
      .Q       (o_data[23]   )
   );

   (* BEL="X13/Y4/lc0" *)
   SB_DFF  dff_2_24 (
      .C       (i_clk         ),
      .D       (p0_dl[25]  ),
      .Q       (p1_dl[24]    )
   );

   (* BEL="X14/Y4/lc0" *)
   SB_DFF  dff_3_24 (
      .C       (i_clk         ),
      .D       (p1_dl[24]    ),
      .Q       (o_data[24]   )
   );

   (* BEL="X13/Y4/lc1" *)
   SB_DFF  dff_2_25 (
      .C       (i_clk         ),
      .D       (p0_dl[26]  ),
      .Q       (p1_dl[25]    )
   );

   (* BEL="X14/Y4/lc1" *)
   SB_DFF  dff_3_25 (
      .C       (i_clk         ),
      .D       (p1_dl[25]    ),
      .Q       (o_data[25]   )
   );

   (* BEL="X13/Y4/lc2" *)
   SB_DFF  dff_2_26 (
      .C       (i_clk         ),
      .D       (p0_dl[27]  ),
      .Q       (p1_dl[26]    )
   );

   (* BEL="X14/Y4/lc2" *)
   SB_DFF  dff_3_26 (
      .C       (i_clk         ),
      .D       (p1_dl[26]    ),
      .Q       (o_data[26]   )
   );

   (* BEL="X13/Y4/lc3" *)
   SB_DFF  dff_2_27 (
      .C       (i_clk         ),
      .D       (p0_dl[28]  ),
      .Q       (p1_dl[27]    )
   );

   (* BEL="X14/Y4/lc3" *)
   SB_DFF  dff_3_27 (
      .C       (i_clk         ),
      .D       (p1_dl[27]    ),
      .Q       (o_data[27]   )
   );

   (* BEL="X13/Y4/lc4" *)
   SB_DFF  dff_2_28 (
      .C       (i_clk         ),
      .D       (p0_dl[29]  ),
      .Q       (p1_dl[28]    )
   );

   (* BEL="X14/Y4/lc4" *)
   SB_DFF  dff_3_28 (
      .C       (i_clk         ),
      .D       (p1_dl[28]    ),
      .Q       (o_data[28]   )
   );

   (* BEL="X13/Y4/lc5" *)
   SB_DFF  dff_2_29 (
      .C       (i_clk         ),
      .D       (p0_dl[30]  ),
      .Q       (p1_dl[29]    )
   );

   (* BEL="X14/Y4/lc5" *)
   SB_DFF  dff_3_29 (
      .C       (i_clk         ),
      .D       (p1_dl[29]    ),
      .Q       (o_data[29]   )
   );

   (* BEL="X13/Y4/lc6" *)
   SB_DFF  dff_2_30 (
      .C       (i_clk         ),
      .D       (p0_dl[31]  ),
      .Q       (p1_dl[30]    )
   );

   (* BEL="X14/Y4/lc6" *)
   SB_DFF  dff_3_30 (
      .C       (i_clk         ),
      .D       (p1_dl[30]    ),
      .Q       (o_data[30]   )
   );

   (* BEL="X13/Y4/lc7" *)
   SB_DFF  dff_2_31 (
      .C       (i_clk         ),
      .D       (p0_dl[32]  ),
      .Q       (p1_dl[31]    )
   );

   (* BEL="X14/Y4/lc7" *)
   SB_DFF  dff_3_31 (
      .C       (i_clk         ),
      .D       (p1_dl[31]    ),
      .Q       (o_data[31]   )
   );

   (* BEL="X13/Y5/lc0" *)
   SB_DFF  dff_2_32 (
      .C       (i_clk         ),
      .D       (p0_dl[33]  ),
      .Q       (p1_dl[32]    )
   );

   (* BEL="X14/Y5/lc0" *)
   SB_DFF  dff_3_32 (
      .C       (i_clk         ),
      .D       (p1_dl[32]    ),
      .Q       (o_data[32]   )
   );

   (* BEL="X13/Y5/lc1" *)
   SB_DFF  dff_2_33 (
      .C       (i_clk         ),
      .D       (p0_dl[34]  ),
      .Q       (p1_dl[33]    )
   );

   (* BEL="X14/Y5/lc1" *)
   SB_DFF  dff_3_33 (
      .C       (i_clk         ),
      .D       (p1_dl[33]    ),
      .Q       (o_data[33]   )
   );

   (* BEL="X13/Y5/lc2" *)
   SB_DFF  dff_2_34 (
      .C       (i_clk         ),
      .D       (p0_dl[35]  ),
      .Q       (p1_dl[34]    )
   );

   (* BEL="X14/Y5/lc2" *)
   SB_DFF  dff_3_34 (
      .C       (i_clk         ),
      .D       (p1_dl[34]    ),
      .Q       (o_data[34]   )
   );

   (* BEL="X13/Y5/lc3" *)
   SB_DFF  dff_2_35 (
      .C       (i_clk         ),
      .D       (p0_dl[36]  ),
      .Q       (p1_dl[35]    )
   );

   (* BEL="X14/Y5/lc3" *)
   SB_DFF  dff_3_35 (
      .C       (i_clk         ),
      .D       (p1_dl[35]    ),
      .Q       (o_data[35]   )
   );

   (* BEL="X13/Y5/lc4" *)
   SB_DFF  dff_2_36 (
      .C       (i_clk         ),
      .D       (p0_dl[37]  ),
      .Q       (p1_dl[36]    )
   );

   (* BEL="X14/Y5/lc4" *)
   SB_DFF  dff_3_36 (
      .C       (i_clk         ),
      .D       (p1_dl[36]    ),
      .Q       (o_data[36]   )
   );

   (* BEL="X13/Y5/lc5" *)
   SB_DFF  dff_2_37 (
      .C       (i_clk         ),
      .D       (p0_dl[38]  ),
      .Q       (p1_dl[37]    )
   );

   (* BEL="X14/Y5/lc5" *)
   SB_DFF  dff_3_37 (
      .C       (i_clk         ),
      .D       (p1_dl[37]    ),
      .Q       (o_data[37]   )
   );

   (* BEL="X13/Y5/lc6" *)
   SB_DFF  dff_2_38 (
      .C       (i_clk         ),
      .D       (p0_dl[39]  ),
      .Q       (p1_dl[38]    )
   );

   (* BEL="X14/Y5/lc6" *)
   SB_DFF  dff_3_38 (
      .C       (i_clk         ),
      .D       (p1_dl[38]    ),
      .Q       (o_data[38]   )
   );

   (* BEL="X13/Y5/lc7" *)
   SB_DFF  dff_2_39 (
      .C       (i_clk         ),
      .D       (p0_dl[40]  ),
      .Q       (p1_dl[39]    )
   );

   (* BEL="X14/Y5/lc7" *)
   SB_DFF  dff_3_39 (
      .C       (i_clk         ),
      .D       (p1_dl[39]    ),
      .Q       (o_data[39]   )
   );

   (* BEL="X13/Y6/lc0" *)
   SB_DFF  dff_2_40 (
      .C       (i_clk         ),
      .D       (p0_dl[41]  ),
      .Q       (p1_dl[40]    )
   );

   (* BEL="X14/Y6/lc0" *)
   SB_DFF  dff_3_40 (
      .C       (i_clk         ),
      .D       (p1_dl[40]    ),
      .Q       (o_data[40]   )
   );

   (* BEL="X13/Y6/lc1" *)
   SB_DFF  dff_2_41 (
      .C       (i_clk         ),
      .D       (p0_dl[42]  ),
      .Q       (p1_dl[41]    )
   );

   (* BEL="X14/Y6/lc1" *)
   SB_DFF  dff_3_41 (
      .C       (i_clk         ),
      .D       (p1_dl[41]    ),
      .Q       (o_data[41]   )
   );

   (* BEL="X13/Y6/lc2" *)
   SB_DFF  dff_2_42 (
      .C       (i_clk         ),
      .D       (p0_dl[43]  ),
      .Q       (p1_dl[42]    )
   );

   (* BEL="X14/Y6/lc2" *)
   SB_DFF  dff_3_42 (
      .C       (i_clk         ),
      .D       (p1_dl[42]    ),
      .Q       (o_data[42]   )
   );

   (* BEL="X13/Y6/lc3" *)
   SB_DFF  dff_2_43 (
      .C       (i_clk         ),
      .D       (p0_dl[44]  ),
      .Q       (p1_dl[43]    )
   );

   (* BEL="X14/Y6/lc3" *)
   SB_DFF  dff_3_43 (
      .C       (i_clk         ),
      .D       (p1_dl[43]    ),
      .Q       (o_data[43]   )
   );

   (* BEL="X13/Y6/lc4" *)
   SB_DFF  dff_2_44 (
      .C       (i_clk         ),
      .D       (p0_dl[45]  ),
      .Q       (p1_dl[44]    )
   );

   (* BEL="X14/Y6/lc4" *)
   SB_DFF  dff_3_44 (
      .C       (i_clk         ),
      .D       (p1_dl[44]    ),
      .Q       (o_data[44]   )
   );

   (* BEL="X13/Y6/lc5" *)
   SB_DFF  dff_2_45 (
      .C       (i_clk         ),
      .D       (p0_dl[46]  ),
      .Q       (p1_dl[45]    )
   );

   (* BEL="X14/Y6/lc5" *)
   SB_DFF  dff_3_45 (
      .C       (i_clk         ),
      .D       (p1_dl[45]    ),
      .Q       (o_data[45]   )
   );

   (* BEL="X13/Y6/lc6" *)
   SB_DFF  dff_2_46 (
      .C       (i_clk         ),
      .D       (p0_dl[47]  ),
      .Q       (p1_dl[46]    )
   );

   (* BEL="X14/Y6/lc6" *)
   SB_DFF  dff_3_46 (
      .C       (i_clk         ),
      .D       (p1_dl[46]    ),
      .Q       (o_data[46]   )
   );

   (* BEL="X13/Y6/lc7" *)
   SB_DFF  dff_2_47 (
      .C       (i_clk         ),
      .D       (p0_dl[48]  ),
      .Q       (p1_dl[47]    )
   );

   (* BEL="X14/Y6/lc7" *)
   SB_DFF  dff_3_47 (
      .C       (i_clk         ),
      .D       (p1_dl[47]    ),
      .Q       (o_data[47]   )
   );

   (* BEL="X13/Y7/lc0" *)
   SB_DFF  dff_2_48 (
      .C       (i_clk         ),
      .D       (p0_dl[49]  ),
      .Q       (p1_dl[48]    )
   );

   (* BEL="X14/Y7/lc0" *)
   SB_DFF  dff_3_48 (
      .C       (i_clk         ),
      .D       (p1_dl[48]    ),
      .Q       (o_data[48]   )
   );

   (* BEL="X13/Y7/lc1" *)
   SB_DFF  dff_2_49 (
      .C       (i_clk         ),
      .D       (p0_dl[50]  ),
      .Q       (p1_dl[49]    )
   );

   (* BEL="X14/Y7/lc1" *)
   SB_DFF  dff_3_49 (
      .C       (i_clk         ),
      .D       (p1_dl[49]    ),
      .Q       (o_data[49]   )
   );

   (* BEL="X13/Y7/lc2" *)
   SB_DFF  dff_2_50 (
      .C       (i_clk         ),
      .D       (p0_dl[51]  ),
      .Q       (p1_dl[50]    )
   );

   (* BEL="X14/Y7/lc2" *)
   SB_DFF  dff_3_50 (
      .C       (i_clk         ),
      .D       (p1_dl[50]    ),
      .Q       (o_data[50]   )
   );

   (* BEL="X13/Y7/lc3" *)
   SB_DFF  dff_2_51 (
      .C       (i_clk         ),
      .D       (p0_dl[52]  ),
      .Q       (p1_dl[51]    )
   );

   (* BEL="X14/Y7/lc3" *)
   SB_DFF  dff_3_51 (
      .C       (i_clk         ),
      .D       (p1_dl[51]    ),
      .Q       (o_data[51]   )
   );

   (* BEL="X13/Y7/lc4" *)
   SB_DFF  dff_2_52 (
      .C       (i_clk         ),
      .D       (p0_dl[53]  ),
      .Q       (p1_dl[52]    )
   );

   (* BEL="X14/Y7/lc4" *)
   SB_DFF  dff_3_52 (
      .C       (i_clk         ),
      .D       (p1_dl[52]    ),
      .Q       (o_data[52]   )
   );

   (* BEL="X13/Y7/lc5" *)
   SB_DFF  dff_2_53 (
      .C       (i_clk         ),
      .D       (p0_dl[54]  ),
      .Q       (p1_dl[53]    )
   );

   (* BEL="X14/Y7/lc5" *)
   SB_DFF  dff_3_53 (
      .C       (i_clk         ),
      .D       (p1_dl[53]    ),
      .Q       (o_data[53]   )
   );

   (* BEL="X13/Y7/lc6" *)
   SB_DFF  dff_2_54 (
      .C       (i_clk         ),
      .D       (p0_dl[55]  ),
      .Q       (p1_dl[54]    )
   );

   (* BEL="X14/Y7/lc6" *)
   SB_DFF  dff_3_54 (
      .C       (i_clk         ),
      .D       (p1_dl[54]    ),
      .Q       (o_data[54]   )
   );

   (* BEL="X13/Y7/lc7" *)
   SB_DFF  dff_2_55 (
      .C       (i_clk         ),
      .D       (p0_dl[56]  ),
      .Q       (p1_dl[55]    )
   );

   (* BEL="X14/Y7/lc7" *)
   SB_DFF  dff_3_55 (
      .C       (i_clk         ),
      .D       (p1_dl[55]    ),
      .Q       (o_data[55]   )
   );

   (* BEL="X13/Y8/lc0" *)
   SB_DFF  dff_2_56 (
      .C       (i_clk         ),
      .D       (p0_dl[57]  ),
      .Q       (p1_dl[56]    )
   );

   (* BEL="X14/Y8/lc0" *)
   SB_DFF  dff_3_56 (
      .C       (i_clk         ),
      .D       (p1_dl[56]    ),
      .Q       (o_data[56]   )
   );

   (* BEL="X13/Y8/lc1" *)
   SB_DFF  dff_2_57 (
      .C       (i_clk         ),
      .D       (p0_dl[58]  ),
      .Q       (p1_dl[57]    )
   );

   (* BEL="X14/Y8/lc1" *)
   SB_DFF  dff_3_57 (
      .C       (i_clk         ),
      .D       (p1_dl[57]    ),
      .Q       (o_data[57]   )
   );

   (* BEL="X13/Y8/lc2" *)
   SB_DFF  dff_2_58 (
      .C       (i_clk         ),
      .D       (p0_dl[59]  ),
      .Q       (p1_dl[58]    )
   );

   (* BEL="X14/Y8/lc2" *)
   SB_DFF  dff_3_58 (
      .C       (i_clk         ),
      .D       (p1_dl[58]    ),
      .Q       (o_data[58]   )
   );

   (* BEL="X13/Y8/lc3" *)
   SB_DFF  dff_2_59 (
      .C       (i_clk         ),
      .D       (p0_dl[60]  ),
      .Q       (p1_dl[59]    )
   );

   (* BEL="X14/Y8/lc3" *)
   SB_DFF  dff_3_59 (
      .C       (i_clk         ),
      .D       (p1_dl[59]    ),
      .Q       (o_data[59]   )
   );

   (* BEL="X13/Y8/lc4" *)
   SB_DFF  dff_2_60 (
      .C       (i_clk         ),
      .D       (p0_dl[61]  ),
      .Q       (p1_dl[60]    )
   );

   (* BEL="X14/Y8/lc4" *)
   SB_DFF  dff_3_60 (
      .C       (i_clk         ),
      .D       (p1_dl[60]    ),
      .Q       (o_data[60]   )
   );

   (* BEL="X13/Y8/lc5" *)
   SB_DFF  dff_2_61 (
      .C       (i_clk         ),
      .D       (p0_dl[62]  ),
      .Q       (p1_dl[61]    )
   );

   (* BEL="X14/Y8/lc5" *)
   SB_DFF  dff_3_61 (
      .C       (i_clk         ),
      .D       (p1_dl[61]    ),
      .Q       (o_data[61]   )
   );

   (* BEL="X13/Y8/lc6" *)
   SB_DFF  dff_2_62 (
      .C       (i_clk         ),
      .D       (p0_dl[63]  ),
      .Q       (p1_dl[62]    )
   );

   (* BEL="X14/Y8/lc6" *)
   SB_DFF  dff_3_62 (
      .C       (i_clk         ),
      .D       (p1_dl[62]    ),
      .Q       (o_data[62]   )
   );

   (* BEL="X13/Y8/lc7" *)
   SB_DFF  dff_2_63 (
      .C       (i_clk         ),
      .D       (p0_dl[64]  ),
      .Q       (p1_dl[63]    )
   );

   (* BEL="X14/Y8/lc7" *)
   SB_DFF  dff_3_63 (
      .C       (i_clk         ),
      .D       (p1_dl[63]    ),
      .Q       (o_data[63]   )
   );

   (* BEL="X13/Y9/lc0" *)
   SB_DFF  dff_2_64 (
      .C       (i_clk         ),
      .D       (p0_dl[65]  ),
      .Q       (p1_dl[64]    )
   );

   (* BEL="X14/Y9/lc0" *)
   SB_DFF  dff_3_64 (
      .C       (i_clk         ),
      .D       (p1_dl[64]    ),
      .Q       (o_data[64]   )
   );

   (* BEL="X13/Y9/lc1" *)
   SB_DFF  dff_2_65 (
      .C       (i_clk         ),
      .D       (p0_dl[66]  ),
      .Q       (p1_dl[65]    )
   );

   (* BEL="X14/Y9/lc1" *)
   SB_DFF  dff_3_65 (
      .C       (i_clk         ),
      .D       (p1_dl[65]    ),
      .Q       (o_data[65]   )
   );

   (* BEL="X13/Y9/lc2" *)
   SB_DFF  dff_2_66 (
      .C       (i_clk         ),
      .D       (p0_dl[67]  ),
      .Q       (p1_dl[66]    )
   );

   (* BEL="X14/Y9/lc2" *)
   SB_DFF  dff_3_66 (
      .C       (i_clk         ),
      .D       (p1_dl[66]    ),
      .Q       (o_data[66]   )
   );

   (* BEL="X13/Y9/lc3" *)
   SB_DFF  dff_2_67 (
      .C       (i_clk         ),
      .D       (p0_dl[68]  ),
      .Q       (p1_dl[67]    )
   );

   (* BEL="X14/Y9/lc3" *)
   SB_DFF  dff_3_67 (
      .C       (i_clk         ),
      .D       (p1_dl[67]    ),
      .Q       (o_data[67]   )
   );

   (* BEL="X13/Y9/lc4" *)
   SB_DFF  dff_2_68 (
      .C       (i_clk         ),
      .D       (p0_dl[69]  ),
      .Q       (p1_dl[68]    )
   );

   (* BEL="X14/Y9/lc4" *)
   SB_DFF  dff_3_68 (
      .C       (i_clk         ),
      .D       (p1_dl[68]    ),
      .Q       (o_data[68]   )
   );

   (* BEL="X13/Y9/lc5" *)
   SB_DFF  dff_2_69 (
      .C       (i_clk         ),
      .D       (p0_dl[70]  ),
      .Q       (p1_dl[69]    )
   );

   (* BEL="X14/Y9/lc5" *)
   SB_DFF  dff_3_69 (
      .C       (i_clk         ),
      .D       (p1_dl[69]    ),
      .Q       (o_data[69]   )
   );

   (* BEL="X13/Y9/lc6" *)
   SB_DFF  dff_2_70 (
      .C       (i_clk         ),
      .D       (p0_dl[71]  ),
      .Q       (p1_dl[70]    )
   );

   (* BEL="X14/Y9/lc6" *)
   SB_DFF  dff_3_70 (
      .C       (i_clk         ),
      .D       (p1_dl[70]    ),
      .Q       (o_data[70]   )
   );

   (* BEL="X13/Y9/lc7" *)
   SB_DFF  dff_2_71 (
      .C       (i_clk         ),
      .D       (p0_dl[72]  ),
      .Q       (p1_dl[71]    )
   );

   (* BEL="X14/Y9/lc7" *)
   SB_DFF  dff_3_71 (
      .C       (i_clk         ),
      .D       (p1_dl[71]    ),
      .Q       (o_data[71]   )
   );

   (* BEL="X13/Y10/lc0" *)
   SB_DFF  dff_2_72 (
      .C       (i_clk         ),
      .D       (p0_dl[73]  ),
      .Q       (p1_dl[72]    )
   );

   (* BEL="X14/Y10/lc0" *)
   SB_DFF  dff_3_72 (
      .C       (i_clk         ),
      .D       (p1_dl[72]    ),
      .Q       (o_data[72]   )
   );

   (* BEL="X13/Y10/lc1" *)
   SB_DFF  dff_2_73 (
      .C       (i_clk         ),
      .D       (p0_dl[74]  ),
      .Q       (p1_dl[73]    )
   );

   (* BEL="X14/Y10/lc1" *)
   SB_DFF  dff_3_73 (
      .C       (i_clk         ),
      .D       (p1_dl[73]    ),
      .Q       (o_data[73]   )
   );

   (* BEL="X13/Y10/lc2" *)
   SB_DFF  dff_2_74 (
      .C       (i_clk         ),
      .D       (p0_dl[75]  ),
      .Q       (p1_dl[74]    )
   );

   (* BEL="X14/Y10/lc2" *)
   SB_DFF  dff_3_74 (
      .C       (i_clk         ),
      .D       (p1_dl[74]    ),
      .Q       (o_data[74]   )
   );

   (* BEL="X13/Y10/lc3" *)
   SB_DFF  dff_2_75 (
      .C       (i_clk         ),
      .D       (p0_dl[76]  ),
      .Q       (p1_dl[75]    )
   );

   (* BEL="X14/Y10/lc3" *)
   SB_DFF  dff_3_75 (
      .C       (i_clk         ),
      .D       (p1_dl[75]    ),
      .Q       (o_data[75]   )
   );

   (* BEL="X13/Y10/lc4" *)
   SB_DFF  dff_2_76 (
      .C       (i_clk         ),
      .D       (p0_dl[77]  ),
      .Q       (p1_dl[76]    )
   );

   (* BEL="X14/Y10/lc4" *)
   SB_DFF  dff_3_76 (
      .C       (i_clk         ),
      .D       (p1_dl[76]    ),
      .Q       (o_data[76]   )
   );

   (* BEL="X13/Y10/lc5" *)
   SB_DFF  dff_2_77 (
      .C       (i_clk         ),
      .D       (p0_dl[78]  ),
      .Q       (p1_dl[77]    )
   );

   (* BEL="X14/Y10/lc5" *)
   SB_DFF  dff_3_77 (
      .C       (i_clk         ),
      .D       (p1_dl[77]    ),
      .Q       (o_data[77]   )
   );

   (* BEL="X13/Y10/lc6" *)
   SB_DFF  dff_2_78 (
      .C       (i_clk         ),
      .D       (p0_dl[79]  ),
      .Q       (p1_dl[78]    )
   );

   (* BEL="X14/Y10/lc6" *)
   SB_DFF  dff_3_78 (
      .C       (i_clk         ),
      .D       (p1_dl[78]    ),
      .Q       (o_data[78]   )
   );

   (* BEL="X13/Y10/lc7" *)
   SB_DFF  dff_2_79 (
      .C       (i_clk         ),
      .D       (p0_dl[80]  ),
      .Q       (p1_dl[79]    )
   );

   (* BEL="X14/Y10/lc7" *)
   SB_DFF  dff_3_79 (
      .C       (i_clk         ),
      .D       (p1_dl[79]    ),
      .Q       (o_data[79]   )
   );

   (* BEL="X13/Y11/lc0" *)
   SB_DFF  dff_2_80 (
      .C       (i_clk         ),
      .D       (p0_dl[81]  ),
      .Q       (p1_dl[80]    )
   );

   (* BEL="X14/Y11/lc0" *)
   SB_DFF  dff_3_80 (
      .C       (i_clk         ),
      .D       (p1_dl[80]    ),
      .Q       (o_data[80]   )
   );

   (* BEL="X13/Y11/lc1" *)
   SB_DFF  dff_2_81 (
      .C       (i_clk         ),
      .D       (p0_dl[82]  ),
      .Q       (p1_dl[81]    )
   );

   (* BEL="X14/Y11/lc1" *)
   SB_DFF  dff_3_81 (
      .C       (i_clk         ),
      .D       (p1_dl[81]    ),
      .Q       (o_data[81]   )
   );

   (* BEL="X13/Y11/lc2" *)
   SB_DFF  dff_2_82 (
      .C       (i_clk         ),
      .D       (p0_dl[83]  ),
      .Q       (p1_dl[82]    )
   );

   (* BEL="X14/Y11/lc2" *)
   SB_DFF  dff_3_82 (
      .C       (i_clk         ),
      .D       (p1_dl[82]    ),
      .Q       (o_data[82]   )
   );

   (* BEL="X13/Y11/lc3" *)
   SB_DFF  dff_2_83 (
      .C       (i_clk         ),
      .D       (p0_dl[84]  ),
      .Q       (p1_dl[83]    )
   );

   (* BEL="X14/Y11/lc3" *)
   SB_DFF  dff_3_83 (
      .C       (i_clk         ),
      .D       (p1_dl[83]    ),
      .Q       (o_data[83]   )
   );

   (* BEL="X13/Y11/lc4" *)
   SB_DFF  dff_2_84 (
      .C       (i_clk         ),
      .D       (p0_dl[85]  ),
      .Q       (p1_dl[84]    )
   );

   (* BEL="X14/Y11/lc4" *)
   SB_DFF  dff_3_84 (
      .C       (i_clk         ),
      .D       (p1_dl[84]    ),
      .Q       (o_data[84]   )
   );

   (* BEL="X13/Y11/lc5" *)
   SB_DFF  dff_2_85 (
      .C       (i_clk         ),
      .D       (p0_dl[86]  ),
      .Q       (p1_dl[85]    )
   );

   (* BEL="X14/Y11/lc5" *)
   SB_DFF  dff_3_85 (
      .C       (i_clk         ),
      .D       (p1_dl[85]    ),
      .Q       (o_data[85]   )
   );

   (* BEL="X13/Y11/lc6" *)
   SB_DFF  dff_2_86 (
      .C       (i_clk         ),
      .D       (p0_dl[87]  ),
      .Q       (p1_dl[86]    )
   );

   (* BEL="X14/Y11/lc6" *)
   SB_DFF  dff_3_86 (
      .C       (i_clk         ),
      .D       (p1_dl[86]    ),
      .Q       (o_data[86]   )
   );

   (* BEL="X13/Y11/lc7" *)
   SB_DFF  dff_2_87 (
      .C       (i_clk         ),
      .D       (p0_dl[88]  ),
      .Q       (p1_dl[87]    )
   );

   (* BEL="X14/Y11/lc7" *)
   SB_DFF  dff_3_87 (
      .C       (i_clk         ),
      .D       (p1_dl[87]    ),
      .Q       (o_data[87]   )
   );

   (* BEL="X13/Y12/lc0" *)
   SB_DFF  dff_2_88 (
      .C       (i_clk         ),
      .D       (p0_dl[89]  ),
      .Q       (p1_dl[88]    )
   );

   (* BEL="X14/Y12/lc0" *)
   SB_DFF  dff_3_88 (
      .C       (i_clk         ),
      .D       (p1_dl[88]    ),
      .Q       (o_data[88]   )
   );

   (* BEL="X13/Y12/lc1" *)
   SB_DFF  dff_2_89 (
      .C       (i_clk         ),
      .D       (p0_dl[90]  ),
      .Q       (p1_dl[89]    )
   );

   (* BEL="X14/Y12/lc1" *)
   SB_DFF  dff_3_89 (
      .C       (i_clk         ),
      .D       (p1_dl[89]    ),
      .Q       (o_data[89]   )
   );

   (* BEL="X13/Y12/lc2" *)
   SB_DFF  dff_2_90 (
      .C       (i_clk         ),
      .D       (p0_dl[91]  ),
      .Q       (p1_dl[90]    )
   );

   (* BEL="X14/Y12/lc2" *)
   SB_DFF  dff_3_90 (
      .C       (i_clk         ),
      .D       (p1_dl[90]    ),
      .Q       (o_data[90]   )
   );

   (* BEL="X13/Y12/lc3" *)
   SB_DFF  dff_2_91 (
      .C       (i_clk         ),
      .D       (p0_dl[92]  ),
      .Q       (p1_dl[91]    )
   );

   (* BEL="X14/Y12/lc3" *)
   SB_DFF  dff_3_91 (
      .C       (i_clk         ),
      .D       (p1_dl[91]    ),
      .Q       (o_data[91]   )
   );

   (* BEL="X13/Y12/lc4" *)
   SB_DFF  dff_2_92 (
      .C       (i_clk         ),
      .D       (p0_dl[93]  ),
      .Q       (p1_dl[92]    )
   );

   (* BEL="X14/Y12/lc4" *)
   SB_DFF  dff_3_92 (
      .C       (i_clk         ),
      .D       (p1_dl[92]    ),
      .Q       (o_data[92]   )
   );

   (* BEL="X13/Y12/lc5" *)
   SB_DFF  dff_2_93 (
      .C       (i_clk         ),
      .D       (p0_dl[94]  ),
      .Q       (p1_dl[93]    )
   );

   (* BEL="X14/Y12/lc5" *)
   SB_DFF  dff_3_93 (
      .C       (i_clk         ),
      .D       (p1_dl[93]    ),
      .Q       (o_data[93]   )
   );

   (* BEL="X13/Y12/lc6" *)
   SB_DFF  dff_2_94 (
      .C       (i_clk         ),
      .D       (p0_dl[95]  ),
      .Q       (p1_dl[94]    )
   );

   (* BEL="X14/Y12/lc6" *)
   SB_DFF  dff_3_94 (
      .C       (i_clk         ),
      .D       (p1_dl[94]    ),
      .Q       (o_data[94]   )
   );

   (* BEL="X13/Y12/lc7" *)
   SB_DFF  dff_2_95 (
      .C       (i_clk         ),
      .D       (p0_dl[96]  ),
      .Q       (p1_dl[95]    )
   );

   (* BEL="X14/Y12/lc7" *)
   SB_DFF  dff_3_95 (
      .C       (i_clk         ),
      .D       (p1_dl[95]    ),
      .Q       (o_data[95]   )
   );

   (* BEL="X13/Y13/lc0" *)
   SB_DFF  dff_2_96 (
      .C       (i_clk         ),
      .D       (p0_dl[97]  ),
      .Q       (p1_dl[96]    )
   );

   (* BEL="X14/Y13/lc0" *)
   SB_DFF  dff_3_96 (
      .C       (i_clk         ),
      .D       (p1_dl[96]    ),
      .Q       (o_data[96]   )
   );

   (* BEL="X13/Y13/lc1" *)
   SB_DFF  dff_2_97 (
      .C       (i_clk         ),
      .D       (p0_dl[98]  ),
      .Q       (p1_dl[97]    )
   );

   (* BEL="X14/Y13/lc1" *)
   SB_DFF  dff_3_97 (
      .C       (i_clk         ),
      .D       (p1_dl[97]    ),
      .Q       (o_data[97]   )
   );

   (* BEL="X13/Y13/lc2" *)
   SB_DFF  dff_2_98 (
      .C       (i_clk         ),
      .D       (p0_dl[99]  ),
      .Q       (p1_dl[98]    )
   );

   (* BEL="X14/Y13/lc2" *)
   SB_DFF  dff_3_98 (
      .C       (i_clk         ),
      .D       (p1_dl[98]    ),
      .Q       (o_data[98]   )
   );

   (* BEL="X13/Y13/lc3" *)
   SB_DFF  dff_2_99 (
      .C       (i_clk         ),
      .D       (p0_dl[100]  ),
      .Q       (p1_dl[99]    )
   );

   (* BEL="X14/Y13/lc3" *)
   SB_DFF  dff_3_99 (
      .C       (i_clk         ),
      .D       (p1_dl[99]    ),
      .Q       (o_data[99]   )
   );

   (* BEL="X13/Y13/lc4" *)
   SB_DFF  dff_2_100 (
      .C       (i_clk         ),
      .D       (p0_dl[101]  ),
      .Q       (p1_dl[100]    )
   );

   (* BEL="X14/Y13/lc4" *)
   SB_DFF  dff_3_100 (
      .C       (i_clk         ),
      .D       (p1_dl[100]    ),
      .Q       (o_data[100]   )
   );

   (* BEL="X13/Y13/lc5" *)
   SB_DFF  dff_2_101 (
      .C       (i_clk         ),
      .D       (p0_dl[102]  ),
      .Q       (p1_dl[101]    )
   );

   (* BEL="X14/Y13/lc5" *)
   SB_DFF  dff_3_101 (
      .C       (i_clk         ),
      .D       (p1_dl[101]    ),
      .Q       (o_data[101]   )
   );

   (* BEL="X13/Y13/lc6" *)
   SB_DFF  dff_2_102 (
      .C       (i_clk         ),
      .D       (p0_dl[103]  ),
      .Q       (p1_dl[102]    )
   );

   (* BEL="X14/Y13/lc6" *)
   SB_DFF  dff_3_102 (
      .C       (i_clk         ),
      .D       (p1_dl[102]    ),
      .Q       (o_data[102]   )
   );

   (* BEL="X13/Y13/lc7" *)
   SB_DFF  dff_2_103 (
      .C       (i_clk         ),
      .D       (p0_dl[104]  ),
      .Q       (p1_dl[103]    )
   );

   (* BEL="X14/Y13/lc7" *)
   SB_DFF  dff_3_103 (
      .C       (i_clk         ),
      .D       (p1_dl[103]    ),
      .Q       (o_data[103]   )
   );

   (* BEL="X13/Y14/lc0" *)
   SB_DFF  dff_2_104 (
      .C       (i_clk         ),
      .D       (p0_dl[105]  ),
      .Q       (p1_dl[104]    )
   );

   (* BEL="X14/Y14/lc0" *)
   SB_DFF  dff_3_104 (
      .C       (i_clk         ),
      .D       (p1_dl[104]    ),
      .Q       (o_data[104]   )
   );

   (* BEL="X13/Y14/lc1" *)
   SB_DFF  dff_2_105 (
      .C       (i_clk         ),
      .D       (p0_dl[106]  ),
      .Q       (p1_dl[105]    )
   );

   (* BEL="X14/Y14/lc1" *)
   SB_DFF  dff_3_105 (
      .C       (i_clk         ),
      .D       (p1_dl[105]    ),
      .Q       (o_data[105]   )
   );

   (* BEL="X13/Y14/lc2" *)
   SB_DFF  dff_2_106 (
      .C       (i_clk         ),
      .D       (p0_dl[107]  ),
      .Q       (p1_dl[106]    )
   );

   (* BEL="X14/Y14/lc2" *)
   SB_DFF  dff_3_106 (
      .C       (i_clk         ),
      .D       (p1_dl[106]    ),
      .Q       (o_data[106]   )
   );

   (* BEL="X13/Y14/lc3" *)
   SB_DFF  dff_2_107 (
      .C       (i_clk         ),
      .D       (p0_dl[108]  ),
      .Q       (p1_dl[107]    )
   );

   (* BEL="X14/Y14/lc3" *)
   SB_DFF  dff_3_107 (
      .C       (i_clk         ),
      .D       (p1_dl[107]    ),
      .Q       (o_data[107]   )
   );

   (* BEL="X13/Y14/lc4" *)
   SB_DFF  dff_2_108 (
      .C       (i_clk         ),
      .D       (p0_dl[109]  ),
      .Q       (p1_dl[108]    )
   );

   (* BEL="X14/Y14/lc4" *)
   SB_DFF  dff_3_108 (
      .C       (i_clk         ),
      .D       (p1_dl[108]    ),
      .Q       (o_data[108]   )
   );

   (* BEL="X13/Y14/lc5" *)
   SB_DFF  dff_2_109 (
      .C       (i_clk         ),
      .D       (p0_dl[110]  ),
      .Q       (p1_dl[109]    )
   );

   (* BEL="X14/Y14/lc5" *)
   SB_DFF  dff_3_109 (
      .C       (i_clk         ),
      .D       (p1_dl[109]    ),
      .Q       (o_data[109]   )
   );

   (* BEL="X13/Y14/lc6" *)
   SB_DFF  dff_2_110 (
      .C       (i_clk         ),
      .D       (p0_dl[111]  ),
      .Q       (p1_dl[110]    )
   );

   (* BEL="X14/Y14/lc6" *)
   SB_DFF  dff_3_110 (
      .C       (i_clk         ),
      .D       (p1_dl[110]    ),
      .Q       (o_data[110]   )
   );

   (* BEL="X13/Y14/lc7" *)
   SB_DFF  dff_2_111 (
      .C       (i_clk         ),
      .D       (p0_dl[112]  ),
      .Q       (p1_dl[111]    )
   );

   (* BEL="X14/Y14/lc7" *)
   SB_DFF  dff_3_111 (
      .C       (i_clk         ),
      .D       (p1_dl[111]    ),
      .Q       (o_data[111]   )
   );

   (* BEL="X13/Y15/lc0" *)
   SB_DFF  dff_2_112 (
      .C       (i_clk         ),
      .D       (p0_dl[113]  ),
      .Q       (p1_dl[112]    )
   );

   (* BEL="X14/Y15/lc0" *)
   SB_DFF  dff_3_112 (
      .C       (i_clk         ),
      .D       (p1_dl[112]    ),
      .Q       (o_data[112]   )
   );

   (* BEL="X13/Y15/lc1" *)
   SB_DFF  dff_2_113 (
      .C       (i_clk         ),
      .D       (p0_dl[114]  ),
      .Q       (p1_dl[113]    )
   );

   (* BEL="X14/Y15/lc1" *)
   SB_DFF  dff_3_113 (
      .C       (i_clk         ),
      .D       (p1_dl[113]    ),
      .Q       (o_data[113]   )
   );

   (* BEL="X13/Y15/lc2" *)
   SB_DFF  dff_2_114 (
      .C       (i_clk         ),
      .D       (p0_dl[115]  ),
      .Q       (p1_dl[114]    )
   );

   (* BEL="X14/Y15/lc2" *)
   SB_DFF  dff_3_114 (
      .C       (i_clk         ),
      .D       (p1_dl[114]    ),
      .Q       (o_data[114]   )
   );

   (* BEL="X13/Y15/lc3" *)
   SB_DFF  dff_2_115 (
      .C       (i_clk         ),
      .D       (p0_dl[116]  ),
      .Q       (p1_dl[115]    )
   );

   (* BEL="X14/Y15/lc3" *)
   SB_DFF  dff_3_115 (
      .C       (i_clk         ),
      .D       (p1_dl[115]    ),
      .Q       (o_data[115]   )
   );

   (* BEL="X13/Y15/lc4" *)
   SB_DFF  dff_2_116 (
      .C       (i_clk         ),
      .D       (p0_dl[117]  ),
      .Q       (p1_dl[116]    )
   );

   (* BEL="X14/Y15/lc4" *)
   SB_DFF  dff_3_116 (
      .C       (i_clk         ),
      .D       (p1_dl[116]    ),
      .Q       (o_data[116]   )
   );

   (* BEL="X13/Y15/lc5" *)
   SB_DFF  dff_2_117 (
      .C       (i_clk         ),
      .D       (p0_dl[118]  ),
      .Q       (p1_dl[117]    )
   );

   (* BEL="X14/Y15/lc5" *)
   SB_DFF  dff_3_117 (
      .C       (i_clk         ),
      .D       (p1_dl[117]    ),
      .Q       (o_data[117]   )
   );

   (* BEL="X13/Y15/lc6" *)
   SB_DFF  dff_2_118 (
      .C       (i_clk         ),
      .D       (p0_dl[119]  ),
      .Q       (p1_dl[118]    )
   );

   (* BEL="X14/Y15/lc6" *)
   SB_DFF  dff_3_118 (
      .C       (i_clk         ),
      .D       (p1_dl[118]    ),
      .Q       (o_data[118]   )
   );

   (* BEL="X13/Y15/lc7" *)
   SB_DFF  dff_2_119 (
      .C       (i_clk         ),
      .D       (p0_dl[120]  ),
      .Q       (p1_dl[119]    )
   );

   (* BEL="X14/Y15/lc7" *)
   SB_DFF  dff_3_119 (
      .C       (i_clk         ),
      .D       (p1_dl[119]    ),
      .Q       (o_data[119]   )
   );

   (* BEL="X13/Y16/lc0" *)
   SB_DFF  dff_2_120 (
      .C       (i_clk         ),
      .D       (p0_dl[121]  ),
      .Q       (p1_dl[120]    )
   );

   (* BEL="X14/Y16/lc0" *)
   SB_DFF  dff_3_120 (
      .C       (i_clk         ),
      .D       (p1_dl[120]    ),
      .Q       (o_data[120]   )
   );

   (* BEL="X13/Y16/lc1" *)
   SB_DFF  dff_2_121 (
      .C       (i_clk         ),
      .D       (p0_dl[122]  ),
      .Q       (p1_dl[121]    )
   );

   (* BEL="X14/Y16/lc1" *)
   SB_DFF  dff_3_121 (
      .C       (i_clk         ),
      .D       (p1_dl[121]    ),
      .Q       (o_data[121]   )
   );

   (* BEL="X13/Y16/lc2" *)
   SB_DFF  dff_2_122 (
      .C       (i_clk         ),
      .D       (p0_dl[123]  ),
      .Q       (p1_dl[122]    )
   );

   (* BEL="X14/Y16/lc2" *)
   SB_DFF  dff_3_122 (
      .C       (i_clk         ),
      .D       (p1_dl[122]    ),
      .Q       (o_data[122]   )
   );

   (* BEL="X13/Y16/lc3" *)
   SB_DFF  dff_2_123 (
      .C       (i_clk         ),
      .D       (p0_dl[124]  ),
      .Q       (p1_dl[123]    )
   );

   (* BEL="X14/Y16/lc3" *)
   SB_DFF  dff_3_123 (
      .C       (i_clk         ),
      .D       (p1_dl[123]    ),
      .Q       (o_data[123]   )
   );

   (* BEL="X13/Y16/lc4" *)
   SB_DFF  dff_2_124 (
      .C       (i_clk         ),
      .D       (p0_dl[125]  ),
      .Q       (p1_dl[124]    )
   );

   (* BEL="X14/Y16/lc4" *)
   SB_DFF  dff_3_124 (
      .C       (i_clk         ),
      .D       (p1_dl[124]    ),
      .Q       (o_data[124]   )
   );

   (* BEL="X13/Y16/lc5" *)
   SB_DFF  dff_2_125 (
      .C       (i_clk         ),
      .D       (p0_dl[126]  ),
      .Q       (p1_dl[125]    )
   );

   (* BEL="X14/Y16/lc5" *)
   SB_DFF  dff_3_125 (
      .C       (i_clk         ),
      .D       (p1_dl[125]    ),
      .Q       (o_data[125]   )
   );

   (* BEL="X13/Y16/lc6" *)
   SB_DFF  dff_2_126 (
      .C       (i_clk         ),
      .D       (p0_dl[127]  ),
      .Q       (p1_dl[126]    )
   );

   (* BEL="X14/Y16/lc6" *)
   SB_DFF  dff_3_126 (
      .C       (i_clk         ),
      .D       (p1_dl[126]    ),
      .Q       (o_data[126]   )
   );

   (* BEL="X13/Y16/lc7" *)
   SB_DFF  dff_2_127 (
      .C       (i_clk         ),
      .D       (p0_dl[128]  ),
      .Q       (p1_dl[127]    )
   );

   (* BEL="X14/Y16/lc7" *)
   SB_DFF  dff_3_127 (
      .C       (i_clk         ),
      .D       (p1_dl[127]    ),
      .Q       (o_data[127]   )
   );

endmodule

